library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity int_to_float is
    port (
        a : in std_logic_vector (23 downto 0);
        b : out std_logic_vector (31 downto 0)
    );
end entity;

architecture rtl of int_to_float is

    -- conversion functions
    function hc_uns(a : std_logic)        return unsigned         is variable b : unsigned(0 downto 0); begin b(0) := a; return b; end;
    function hc_uns(a : std_logic_vector) return unsigned         is begin return unsigned(a); end;
    function hc_sgn(a : std_logic)        return signed           is variable b : signed(0 downto 0); begin b(0) := a; return b; end;
    function hc_sgn(a : std_logic_vector) return signed           is begin return signed(a); end;
    function hc_sl (a : std_logic_vector) return std_logic        is begin return a(a'right); end;
    function hc_sl (a : unsigned)         return std_logic        is begin return a(a'right); end;
    function hc_sl (a : signed)           return std_logic        is begin return a(a'right); end;
    function hc_sl (a : boolean)          return std_logic        is begin if a then return '1'; else return '0'; end if; end;
    function hc_slv(a : std_logic_vector) return std_logic_vector is begin return a; end;
    function hc_slv(a : unsigned)         return std_logic_vector is begin return std_logic_vector(a); end;
    function hc_slv(a : signed)           return std_logic_vector is begin return std_logic_vector(a); end;

    -- signal declarations
    constant hc_935 : std_logic_vector (31 downto 0) := "00000000000000000000000000000000";
    signal hc_933 : std_logic;
    signal hc_932 : std_logic;
    signal hc_931 : std_logic;
    signal hc_930 : std_logic;
    signal hc_929 : std_logic;
    signal hc_928 : std_logic;
    signal hc_927 : std_logic;
    signal hc_926 : std_logic;
    signal hc_925 : std_logic;
    signal hc_924 : std_logic;
    signal hc_923 : std_logic;
    signal hc_922 : std_logic;
    signal hc_921 : std_logic;
    signal hc_920 : std_logic;
    signal hc_919 : std_logic;
    signal hc_918 : std_logic;
    signal hc_917 : std_logic;
    signal hc_916 : std_logic;
    signal hc_915 : std_logic;
    signal hc_914 : std_logic;
    signal hc_913 : std_logic;
    signal hc_912 : std_logic;
    signal hc_903 : std_logic;
    signal hc_902 : std_logic;
    signal hc_901 : std_logic;
    signal hc_900 : std_logic;
    signal hc_899 : std_logic;
    signal hc_898 : std_logic;
    signal hc_897 : std_logic;
    signal hc_896 : std_logic;
    signal hc_895 : std_logic;
    signal hc_894 : std_logic;
    signal hc_893 : std_logic;
    signal hc_892 : std_logic;
    signal hc_891 : std_logic;
    signal hc_890 : std_logic;
    signal hc_889 : std_logic;
    signal hc_888 : std_logic;
    signal hc_887 : std_logic;
    signal hc_886 : std_logic;
    signal hc_885 : std_logic;
    signal hc_884 : std_logic;
    signal hc_883 : std_logic;
    signal hc_882 : std_logic;
    constant hc_879 : std_logic := '0';
    signal hc_878 : std_logic_vector (22 downto 0);
    signal hc_880 : std_logic_vector (23 downto 0);
    signal hc_881 : std_logic;
    signal hc_904 : std_logic_vector (22 downto 0);
    signal hc_876 : std_logic;
    signal hc_875 : std_logic;
    signal hc_874 : std_logic;
    signal hc_873 : std_logic;
    signal hc_872 : std_logic;
    signal hc_871 : std_logic;
    signal hc_870 : std_logic;
    signal hc_869 : std_logic;
    signal hc_868 : std_logic;
    signal hc_867 : std_logic;
    signal hc_866 : std_logic;
    signal hc_865 : std_logic;
    signal hc_864 : std_logic;
    signal hc_863 : std_logic;
    signal hc_862 : std_logic;
    signal hc_861 : std_logic;
    signal hc_860 : std_logic;
    signal hc_859 : std_logic;
    signal hc_858 : std_logic;
    signal hc_857 : std_logic;
    signal hc_856 : std_logic;
    signal hc_855 : std_logic;
    constant hc_852 : std_logic_vector (1 downto 0) := "00";
    signal hc_851 : std_logic_vector (21 downto 0);
    signal hc_853 : std_logic_vector (23 downto 0);
    signal hc_854 : std_logic;
    signal hc_877 : std_logic_vector (22 downto 0);
    signal hc_905 : std_logic_vector (22 downto 0);
    signal hc_848 : std_logic;
    signal hc_847 : std_logic;
    signal hc_846 : std_logic;
    signal hc_845 : std_logic;
    signal hc_844 : std_logic;
    signal hc_843 : std_logic;
    signal hc_842 : std_logic;
    signal hc_841 : std_logic;
    signal hc_840 : std_logic;
    signal hc_839 : std_logic;
    signal hc_838 : std_logic;
    signal hc_837 : std_logic;
    signal hc_836 : std_logic;
    signal hc_835 : std_logic;
    signal hc_834 : std_logic;
    signal hc_833 : std_logic;
    signal hc_832 : std_logic;
    signal hc_831 : std_logic;
    signal hc_830 : std_logic;
    signal hc_829 : std_logic;
    signal hc_828 : std_logic;
    signal hc_827 : std_logic;
    constant hc_824 : std_logic_vector (2 downto 0) := "000";
    signal hc_823 : std_logic_vector (20 downto 0);
    signal hc_825 : std_logic_vector (23 downto 0);
    signal hc_826 : std_logic;
    signal hc_849 : std_logic_vector (22 downto 0);
    signal hc_821 : std_logic;
    signal hc_820 : std_logic;
    signal hc_819 : std_logic;
    signal hc_818 : std_logic;
    signal hc_817 : std_logic;
    signal hc_816 : std_logic;
    signal hc_815 : std_logic;
    signal hc_814 : std_logic;
    signal hc_813 : std_logic;
    signal hc_812 : std_logic;
    signal hc_811 : std_logic;
    signal hc_810 : std_logic;
    signal hc_809 : std_logic;
    signal hc_808 : std_logic;
    signal hc_807 : std_logic;
    signal hc_806 : std_logic;
    signal hc_805 : std_logic;
    signal hc_804 : std_logic;
    signal hc_803 : std_logic;
    signal hc_802 : std_logic;
    signal hc_801 : std_logic;
    signal hc_800 : std_logic;
    constant hc_797 : std_logic_vector (3 downto 0) := "0000";
    signal hc_796 : std_logic_vector (19 downto 0);
    signal hc_798 : std_logic_vector (23 downto 0);
    signal hc_799 : std_logic;
    signal hc_822 : std_logic_vector (22 downto 0);
    signal hc_850 : std_logic_vector (22 downto 0);
    signal hc_906 : std_logic_vector (22 downto 0);
    signal hc_792 : std_logic;
    signal hc_791 : std_logic;
    signal hc_790 : std_logic;
    signal hc_789 : std_logic;
    signal hc_788 : std_logic;
    signal hc_787 : std_logic;
    signal hc_786 : std_logic;
    signal hc_785 : std_logic;
    signal hc_784 : std_logic;
    signal hc_783 : std_logic;
    signal hc_782 : std_logic;
    signal hc_781 : std_logic;
    signal hc_780 : std_logic;
    signal hc_779 : std_logic;
    signal hc_778 : std_logic;
    signal hc_777 : std_logic;
    signal hc_776 : std_logic;
    signal hc_775 : std_logic;
    signal hc_774 : std_logic;
    signal hc_773 : std_logic;
    signal hc_772 : std_logic;
    signal hc_771 : std_logic;
    constant hc_768 : std_logic_vector (4 downto 0) := "00000";
    signal hc_767 : std_logic_vector (18 downto 0);
    signal hc_769 : std_logic_vector (23 downto 0);
    signal hc_770 : std_logic;
    signal hc_793 : std_logic_vector (22 downto 0);
    signal hc_765 : std_logic;
    signal hc_764 : std_logic;
    signal hc_763 : std_logic;
    signal hc_762 : std_logic;
    signal hc_761 : std_logic;
    signal hc_760 : std_logic;
    signal hc_759 : std_logic;
    signal hc_758 : std_logic;
    signal hc_757 : std_logic;
    signal hc_756 : std_logic;
    signal hc_755 : std_logic;
    signal hc_754 : std_logic;
    signal hc_753 : std_logic;
    signal hc_752 : std_logic;
    signal hc_751 : std_logic;
    signal hc_750 : std_logic;
    signal hc_749 : std_logic;
    signal hc_748 : std_logic;
    signal hc_747 : std_logic;
    signal hc_746 : std_logic;
    signal hc_745 : std_logic;
    signal hc_744 : std_logic;
    constant hc_741 : std_logic_vector (5 downto 0) := "000000";
    signal hc_740 : std_logic_vector (17 downto 0);
    signal hc_742 : std_logic_vector (23 downto 0);
    signal hc_743 : std_logic;
    signal hc_766 : std_logic_vector (22 downto 0);
    signal hc_794 : std_logic_vector (22 downto 0);
    signal hc_737 : std_logic;
    signal hc_736 : std_logic;
    signal hc_735 : std_logic;
    signal hc_734 : std_logic;
    signal hc_733 : std_logic;
    signal hc_732 : std_logic;
    signal hc_731 : std_logic;
    signal hc_730 : std_logic;
    signal hc_729 : std_logic;
    signal hc_728 : std_logic;
    signal hc_727 : std_logic;
    signal hc_726 : std_logic;
    signal hc_725 : std_logic;
    signal hc_724 : std_logic;
    signal hc_723 : std_logic;
    signal hc_722 : std_logic;
    signal hc_721 : std_logic;
    signal hc_720 : std_logic;
    signal hc_719 : std_logic;
    signal hc_718 : std_logic;
    signal hc_717 : std_logic;
    signal hc_716 : std_logic;
    constant hc_713 : std_logic_vector (6 downto 0) := "0000000";
    signal hc_712 : std_logic_vector (16 downto 0);
    signal hc_714 : std_logic_vector (23 downto 0);
    signal hc_715 : std_logic;
    signal hc_738 : std_logic_vector (22 downto 0);
    signal hc_710 : std_logic;
    signal hc_709 : std_logic;
    signal hc_708 : std_logic;
    signal hc_707 : std_logic;
    signal hc_706 : std_logic;
    signal hc_705 : std_logic;
    signal hc_704 : std_logic;
    signal hc_703 : std_logic;
    signal hc_702 : std_logic;
    signal hc_701 : std_logic;
    signal hc_700 : std_logic;
    signal hc_699 : std_logic;
    signal hc_698 : std_logic;
    signal hc_697 : std_logic;
    signal hc_696 : std_logic;
    signal hc_695 : std_logic;
    signal hc_694 : std_logic;
    signal hc_693 : std_logic;
    signal hc_692 : std_logic;
    signal hc_691 : std_logic;
    signal hc_690 : std_logic;
    signal hc_689 : std_logic;
    constant hc_686 : std_logic_vector (7 downto 0) := "00000000";
    signal hc_685 : std_logic_vector (15 downto 0);
    signal hc_687 : std_logic_vector (23 downto 0);
    signal hc_688 : std_logic;
    signal hc_711 : std_logic_vector (22 downto 0);
    signal hc_739 : std_logic_vector (22 downto 0);
    signal hc_795 : std_logic_vector (22 downto 0);
    signal hc_907 : std_logic_vector (22 downto 0);
    signal hc_680 : std_logic;
    signal hc_679 : std_logic;
    signal hc_678 : std_logic;
    signal hc_677 : std_logic;
    signal hc_676 : std_logic;
    signal hc_675 : std_logic;
    signal hc_674 : std_logic;
    signal hc_673 : std_logic;
    signal hc_672 : std_logic;
    signal hc_671 : std_logic;
    signal hc_670 : std_logic;
    signal hc_669 : std_logic;
    signal hc_668 : std_logic;
    signal hc_667 : std_logic;
    signal hc_666 : std_logic;
    signal hc_665 : std_logic;
    signal hc_664 : std_logic;
    signal hc_663 : std_logic;
    signal hc_662 : std_logic;
    signal hc_661 : std_logic;
    signal hc_660 : std_logic;
    signal hc_659 : std_logic;
    constant hc_656 : std_logic_vector (8 downto 0) := "000000000";
    signal hc_655 : std_logic_vector (14 downto 0);
    signal hc_657 : std_logic_vector (23 downto 0);
    signal hc_658 : std_logic;
    signal hc_681 : std_logic_vector (22 downto 0);
    signal hc_653 : std_logic;
    signal hc_652 : std_logic;
    signal hc_651 : std_logic;
    signal hc_650 : std_logic;
    signal hc_649 : std_logic;
    signal hc_648 : std_logic;
    signal hc_647 : std_logic;
    signal hc_646 : std_logic;
    signal hc_645 : std_logic;
    signal hc_644 : std_logic;
    signal hc_643 : std_logic;
    signal hc_642 : std_logic;
    signal hc_641 : std_logic;
    signal hc_640 : std_logic;
    signal hc_639 : std_logic;
    signal hc_638 : std_logic;
    signal hc_637 : std_logic;
    signal hc_636 : std_logic;
    signal hc_635 : std_logic;
    signal hc_634 : std_logic;
    signal hc_633 : std_logic;
    signal hc_632 : std_logic;
    constant hc_629 : std_logic_vector (9 downto 0) := "0000000000";
    signal hc_628 : std_logic_vector (13 downto 0);
    signal hc_630 : std_logic_vector (23 downto 0);
    signal hc_631 : std_logic;
    signal hc_654 : std_logic_vector (22 downto 0);
    signal hc_682 : std_logic_vector (22 downto 0);
    signal hc_625 : std_logic;
    signal hc_624 : std_logic;
    signal hc_623 : std_logic;
    signal hc_622 : std_logic;
    signal hc_621 : std_logic;
    signal hc_620 : std_logic;
    signal hc_619 : std_logic;
    signal hc_618 : std_logic;
    signal hc_617 : std_logic;
    signal hc_616 : std_logic;
    signal hc_615 : std_logic;
    signal hc_614 : std_logic;
    signal hc_613 : std_logic;
    signal hc_612 : std_logic;
    signal hc_611 : std_logic;
    signal hc_610 : std_logic;
    signal hc_609 : std_logic;
    signal hc_608 : std_logic;
    signal hc_607 : std_logic;
    signal hc_606 : std_logic;
    signal hc_605 : std_logic;
    signal hc_604 : std_logic;
    constant hc_601 : std_logic_vector (10 downto 0) := "00000000000";
    signal hc_600 : std_logic_vector (12 downto 0);
    signal hc_602 : std_logic_vector (23 downto 0);
    signal hc_603 : std_logic;
    signal hc_626 : std_logic_vector (22 downto 0);
    signal hc_598 : std_logic;
    signal hc_597 : std_logic;
    signal hc_596 : std_logic;
    signal hc_595 : std_logic;
    signal hc_594 : std_logic;
    signal hc_593 : std_logic;
    signal hc_592 : std_logic;
    signal hc_591 : std_logic;
    signal hc_590 : std_logic;
    signal hc_589 : std_logic;
    signal hc_588 : std_logic;
    signal hc_587 : std_logic;
    signal hc_586 : std_logic;
    signal hc_585 : std_logic;
    signal hc_584 : std_logic;
    signal hc_583 : std_logic;
    signal hc_582 : std_logic;
    signal hc_581 : std_logic;
    signal hc_580 : std_logic;
    signal hc_579 : std_logic;
    signal hc_578 : std_logic;
    signal hc_577 : std_logic;
    constant hc_574 : std_logic_vector (11 downto 0) := "000000000000";
    signal hc_573 : std_logic_vector (11 downto 0);
    signal hc_575 : std_logic_vector (23 downto 0);
    signal hc_576 : std_logic;
    signal hc_599 : std_logic_vector (22 downto 0);
    signal hc_627 : std_logic_vector (22 downto 0);
    signal hc_683 : std_logic_vector (22 downto 0);
    signal hc_569 : std_logic;
    signal hc_568 : std_logic;
    signal hc_567 : std_logic;
    signal hc_566 : std_logic;
    signal hc_565 : std_logic;
    signal hc_564 : std_logic;
    signal hc_563 : std_logic;
    signal hc_562 : std_logic;
    signal hc_561 : std_logic;
    signal hc_560 : std_logic;
    signal hc_559 : std_logic;
    signal hc_558 : std_logic;
    signal hc_557 : std_logic;
    signal hc_556 : std_logic;
    signal hc_555 : std_logic;
    signal hc_554 : std_logic;
    signal hc_553 : std_logic;
    signal hc_552 : std_logic;
    signal hc_551 : std_logic;
    signal hc_550 : std_logic;
    signal hc_549 : std_logic;
    signal hc_548 : std_logic;
    constant hc_545 : std_logic_vector (12 downto 0) := "0000000000000";
    signal hc_544 : std_logic_vector (10 downto 0);
    signal hc_546 : std_logic_vector (23 downto 0);
    signal hc_547 : std_logic;
    signal hc_570 : std_logic_vector (22 downto 0);
    signal hc_542 : std_logic;
    signal hc_541 : std_logic;
    signal hc_540 : std_logic;
    signal hc_539 : std_logic;
    signal hc_538 : std_logic;
    signal hc_537 : std_logic;
    signal hc_536 : std_logic;
    signal hc_535 : std_logic;
    signal hc_534 : std_logic;
    signal hc_533 : std_logic;
    signal hc_532 : std_logic;
    signal hc_531 : std_logic;
    signal hc_530 : std_logic;
    signal hc_529 : std_logic;
    signal hc_528 : std_logic;
    signal hc_527 : std_logic;
    signal hc_526 : std_logic;
    signal hc_525 : std_logic;
    signal hc_524 : std_logic;
    signal hc_523 : std_logic;
    signal hc_522 : std_logic;
    signal hc_521 : std_logic;
    constant hc_518 : std_logic_vector (13 downto 0) := "00000000000000";
    signal hc_517 : std_logic_vector (9 downto 0);
    signal hc_519 : std_logic_vector (23 downto 0);
    signal hc_520 : std_logic;
    signal hc_543 : std_logic_vector (22 downto 0);
    signal hc_571 : std_logic_vector (22 downto 0);
    signal hc_514 : std_logic;
    signal hc_513 : std_logic;
    signal hc_512 : std_logic;
    signal hc_511 : std_logic;
    signal hc_510 : std_logic;
    signal hc_509 : std_logic;
    signal hc_508 : std_logic;
    signal hc_507 : std_logic;
    signal hc_506 : std_logic;
    signal hc_505 : std_logic;
    signal hc_504 : std_logic;
    signal hc_503 : std_logic;
    signal hc_502 : std_logic;
    signal hc_501 : std_logic;
    signal hc_500 : std_logic;
    signal hc_499 : std_logic;
    signal hc_498 : std_logic;
    signal hc_497 : std_logic;
    signal hc_496 : std_logic;
    signal hc_495 : std_logic;
    signal hc_494 : std_logic;
    signal hc_493 : std_logic;
    constant hc_490 : std_logic_vector (14 downto 0) := "000000000000000";
    signal hc_489 : std_logic_vector (8 downto 0);
    signal hc_491 : std_logic_vector (23 downto 0);
    signal hc_492 : std_logic;
    signal hc_515 : std_logic_vector (22 downto 0);
    signal hc_487 : std_logic;
    signal hc_486 : std_logic;
    signal hc_485 : std_logic;
    signal hc_484 : std_logic;
    signal hc_483 : std_logic;
    signal hc_482 : std_logic;
    signal hc_481 : std_logic;
    signal hc_480 : std_logic;
    signal hc_479 : std_logic;
    signal hc_478 : std_logic;
    signal hc_477 : std_logic;
    signal hc_476 : std_logic;
    signal hc_475 : std_logic;
    signal hc_474 : std_logic;
    signal hc_473 : std_logic;
    signal hc_472 : std_logic;
    signal hc_471 : std_logic;
    signal hc_470 : std_logic;
    signal hc_469 : std_logic;
    signal hc_468 : std_logic;
    signal hc_467 : std_logic;
    signal hc_466 : std_logic;
    constant hc_463 : std_logic_vector (15 downto 0) := "0000000000000000";
    signal hc_462 : std_logic_vector (7 downto 0);
    signal hc_464 : std_logic_vector (23 downto 0);
    signal hc_465 : std_logic;
    signal hc_488 : std_logic_vector (22 downto 0);
    signal hc_516 : std_logic_vector (22 downto 0);
    signal hc_572 : std_logic_vector (22 downto 0);
    signal hc_684 : std_logic_vector (22 downto 0);
    signal hc_908 : std_logic_vector (22 downto 0);
    signal hc_457 : std_logic;
    signal hc_456 : std_logic;
    signal hc_455 : std_logic;
    signal hc_454 : std_logic;
    signal hc_453 : std_logic;
    signal hc_452 : std_logic;
    signal hc_451 : std_logic;
    signal hc_450 : std_logic;
    signal hc_449 : std_logic;
    signal hc_448 : std_logic;
    signal hc_447 : std_logic;
    signal hc_446 : std_logic;
    signal hc_445 : std_logic;
    signal hc_444 : std_logic;
    signal hc_443 : std_logic;
    signal hc_442 : std_logic;
    signal hc_441 : std_logic;
    signal hc_440 : std_logic;
    signal hc_439 : std_logic;
    signal hc_438 : std_logic;
    signal hc_437 : std_logic;
    signal hc_436 : std_logic;
    constant hc_433 : std_logic_vector (16 downto 0) := "00000000000000000";
    signal hc_432 : std_logic_vector (6 downto 0);
    signal hc_434 : std_logic_vector (23 downto 0);
    signal hc_435 : std_logic;
    signal hc_458 : std_logic_vector (22 downto 0);
    signal hc_430 : std_logic;
    signal hc_429 : std_logic;
    signal hc_428 : std_logic;
    signal hc_427 : std_logic;
    signal hc_426 : std_logic;
    signal hc_425 : std_logic;
    signal hc_424 : std_logic;
    signal hc_423 : std_logic;
    signal hc_422 : std_logic;
    signal hc_421 : std_logic;
    signal hc_420 : std_logic;
    signal hc_419 : std_logic;
    signal hc_418 : std_logic;
    signal hc_417 : std_logic;
    signal hc_416 : std_logic;
    signal hc_415 : std_logic;
    signal hc_414 : std_logic;
    signal hc_413 : std_logic;
    signal hc_412 : std_logic;
    signal hc_411 : std_logic;
    signal hc_410 : std_logic;
    signal hc_409 : std_logic;
    constant hc_406 : std_logic_vector (17 downto 0) := "000000000000000000";
    signal hc_405 : std_logic_vector (5 downto 0);
    signal hc_407 : std_logic_vector (23 downto 0);
    signal hc_408 : std_logic;
    signal hc_431 : std_logic_vector (22 downto 0);
    signal hc_459 : std_logic_vector (22 downto 0);
    signal hc_402 : std_logic;
    signal hc_401 : std_logic;
    signal hc_400 : std_logic;
    signal hc_399 : std_logic;
    signal hc_398 : std_logic;
    signal hc_397 : std_logic;
    signal hc_396 : std_logic;
    signal hc_395 : std_logic;
    signal hc_394 : std_logic;
    signal hc_393 : std_logic;
    signal hc_392 : std_logic;
    signal hc_391 : std_logic;
    signal hc_390 : std_logic;
    signal hc_389 : std_logic;
    signal hc_388 : std_logic;
    signal hc_387 : std_logic;
    signal hc_386 : std_logic;
    signal hc_385 : std_logic;
    signal hc_384 : std_logic;
    signal hc_383 : std_logic;
    signal hc_382 : std_logic;
    signal hc_381 : std_logic;
    constant hc_378 : std_logic_vector (18 downto 0) := "0000000000000000000";
    signal hc_377 : std_logic_vector (4 downto 0);
    signal hc_379 : std_logic_vector (23 downto 0);
    signal hc_380 : std_logic;
    signal hc_403 : std_logic_vector (22 downto 0);
    signal hc_375 : std_logic;
    signal hc_374 : std_logic;
    signal hc_373 : std_logic;
    signal hc_372 : std_logic;
    signal hc_371 : std_logic;
    signal hc_370 : std_logic;
    signal hc_369 : std_logic;
    signal hc_368 : std_logic;
    signal hc_367 : std_logic;
    signal hc_366 : std_logic;
    signal hc_365 : std_logic;
    signal hc_364 : std_logic;
    signal hc_363 : std_logic;
    signal hc_362 : std_logic;
    signal hc_361 : std_logic;
    signal hc_360 : std_logic;
    signal hc_359 : std_logic;
    signal hc_358 : std_logic;
    signal hc_357 : std_logic;
    signal hc_356 : std_logic;
    signal hc_355 : std_logic;
    signal hc_354 : std_logic;
    constant hc_351 : std_logic_vector (19 downto 0) := "00000000000000000000";
    signal hc_350 : std_logic_vector (3 downto 0);
    signal hc_352 : std_logic_vector (23 downto 0);
    signal hc_353 : std_logic;
    signal hc_376 : std_logic_vector (22 downto 0);
    signal hc_404 : std_logic_vector (22 downto 0);
    signal hc_460 : std_logic_vector (22 downto 0);
    signal hc_346 : std_logic;
    signal hc_345 : std_logic;
    signal hc_344 : std_logic;
    signal hc_343 : std_logic;
    signal hc_342 : std_logic;
    signal hc_341 : std_logic;
    signal hc_340 : std_logic;
    signal hc_339 : std_logic;
    signal hc_338 : std_logic;
    signal hc_337 : std_logic;
    signal hc_336 : std_logic;
    signal hc_335 : std_logic;
    signal hc_334 : std_logic;
    signal hc_333 : std_logic;
    signal hc_332 : std_logic;
    signal hc_331 : std_logic;
    signal hc_330 : std_logic;
    signal hc_329 : std_logic;
    signal hc_328 : std_logic;
    signal hc_327 : std_logic;
    signal hc_326 : std_logic;
    signal hc_325 : std_logic;
    constant hc_322 : std_logic_vector (20 downto 0) := "000000000000000000000";
    signal hc_321 : std_logic_vector (2 downto 0);
    signal hc_323 : std_logic_vector (23 downto 0);
    signal hc_324 : std_logic;
    signal hc_347 : std_logic_vector (22 downto 0);
    signal hc_319 : std_logic;
    signal hc_318 : std_logic;
    signal hc_317 : std_logic;
    signal hc_316 : std_logic;
    signal hc_315 : std_logic;
    signal hc_314 : std_logic;
    signal hc_313 : std_logic;
    signal hc_312 : std_logic;
    signal hc_311 : std_logic;
    signal hc_310 : std_logic;
    signal hc_309 : std_logic;
    signal hc_308 : std_logic;
    signal hc_307 : std_logic;
    signal hc_306 : std_logic;
    signal hc_305 : std_logic;
    signal hc_304 : std_logic;
    signal hc_303 : std_logic;
    signal hc_302 : std_logic;
    signal hc_301 : std_logic;
    signal hc_300 : std_logic;
    signal hc_299 : std_logic;
    signal hc_298 : std_logic;
    constant hc_295 : std_logic_vector (21 downto 0) := "0000000000000000000000";
    signal hc_294 : std_logic_vector (1 downto 0);
    signal hc_296 : std_logic_vector (23 downto 0);
    signal hc_297 : std_logic;
    signal hc_320 : std_logic_vector (22 downto 0);
    signal hc_348 : std_logic_vector (22 downto 0);
    signal hc_291 : std_logic;
    signal hc_290 : std_logic;
    signal hc_289 : std_logic;
    signal hc_288 : std_logic;
    signal hc_287 : std_logic;
    signal hc_286 : std_logic;
    signal hc_285 : std_logic;
    signal hc_284 : std_logic;
    signal hc_283 : std_logic;
    signal hc_282 : std_logic;
    signal hc_281 : std_logic;
    signal hc_280 : std_logic;
    signal hc_279 : std_logic;
    signal hc_278 : std_logic;
    signal hc_277 : std_logic;
    signal hc_276 : std_logic;
    signal hc_275 : std_logic;
    signal hc_274 : std_logic;
    signal hc_273 : std_logic;
    signal hc_272 : std_logic;
    signal hc_271 : std_logic;
    signal hc_270 : std_logic;
    constant hc_267 : std_logic_vector (22 downto 0) := "00000000000000000000000";
    signal hc_266 : std_logic;
    signal hc_268 : std_logic_vector (23 downto 0);
    signal hc_269 : std_logic;
    signal hc_292 : std_logic_vector (22 downto 0);
    constant hc_265 : std_logic_vector (22 downto 0) := "00000000000000000000000";
    signal hc_293 : std_logic_vector (22 downto 0);
    signal hc_349 : std_logic_vector (22 downto 0);
    signal hc_461 : std_logic_vector (22 downto 0);
    signal hc_909 : std_logic_vector (22 downto 0);
    constant hc_264 : std_logic_vector (22 downto 0) := "00000000000000000000000";
    signal hc_259 : std_logic;
    signal hc_258 : std_logic;
    signal hc_260 : std_logic;
    signal hc_256 : std_logic;
    signal hc_255 : std_logic;
    signal hc_257 : std_logic;
    signal hc_261 : std_logic;
    signal hc_252 : std_logic;
    signal hc_251 : std_logic;
    signal hc_253 : std_logic;
    signal hc_249 : std_logic;
    signal hc_248 : std_logic;
    signal hc_250 : std_logic;
    signal hc_254 : std_logic;
    signal hc_262 : std_logic;
    signal hc_243 : std_logic;
    signal hc_242 : std_logic;
    signal hc_244 : std_logic;
    signal hc_240 : std_logic;
    signal hc_239 : std_logic;
    signal hc_241 : std_logic;
    signal hc_245 : std_logic;
    signal hc_236 : std_logic;
    signal hc_235 : std_logic;
    signal hc_237 : std_logic;
    signal hc_233 : std_logic;
    signal hc_232 : std_logic;
    signal hc_234 : std_logic;
    signal hc_238 : std_logic;
    signal hc_246 : std_logic;
    signal hc_228 : std_logic;
    signal hc_227 : std_logic;
    signal hc_229 : std_logic;
    signal hc_225 : std_logic;
    signal hc_224 : std_logic;
    signal hc_226 : std_logic;
    signal hc_230 : std_logic;
    signal hc_221 : std_logic;
    signal hc_220 : std_logic;
    signal hc_222 : std_logic;
    signal hc_218 : std_logic;
    signal hc_215 : std_logic;
    signal hc_214 : std_logic;
    signal hc_213 : std_logic;
    signal hc_212 : std_logic;
    signal hc_211 : std_logic;
    signal hc_210 : std_logic;
    signal hc_209 : std_logic;
    signal hc_208 : std_logic;
    signal hc_207 : std_logic;
    signal hc_206 : std_logic;
    signal hc_205 : std_logic;
    signal hc_204 : std_logic;
    signal hc_203 : std_logic;
    signal hc_202 : std_logic;
    signal hc_201 : std_logic;
    signal hc_200 : std_logic;
    signal hc_199 : std_logic;
    signal hc_198 : std_logic;
    signal hc_197 : std_logic;
    signal hc_196 : std_logic;
    signal hc_195 : std_logic;
    signal hc_194 : std_logic;
    signal hc_193 : std_logic;
    signal hc_192 : std_logic;
    signal hc_216 : std_logic_vector (23 downto 0);
    signal hc_217 : std_logic;
    signal hc_219 : std_logic;
    signal hc_223 : std_logic;
    signal hc_231 : std_logic;
    signal hc_247 : std_logic;
    signal hc_263 : std_logic;
    signal hc_910 : std_logic_vector (22 downto 0);
    signal hc_911 : std_logic;
    signal hc_191 : std_logic;
    signal hc_190 : std_logic;
    signal hc_189 : std_logic;
    signal hc_188 : std_logic;
    signal hc_187 : std_logic;
    signal hc_186 : std_logic;
    signal hc_185 : std_logic;
    constant hc_182 : std_logic_vector (7 downto 0) := "01111111";
    constant hc_180 : std_logic_vector (7 downto 0) := "00000001";
    signal hc_181 : std_logic_vector (7 downto 0);
    signal hc_183 : std_logic_vector (7 downto 0);
    signal hc_184 : std_logic;
    signal hc_179 : std_logic;
    signal hc_934 : std_logic_vector (31 downto 0);
    constant hc_177 : std_logic_vector (7 downto 0) := "00000000";
    constant hc_170 : std_logic_vector (7 downto 0) := "00011000";
    constant hc_169 : std_logic_vector (7 downto 0) := "00010111";
    signal hc_171 : std_logic_vector (7 downto 0);
    constant hc_167 : std_logic_vector (7 downto 0) := "00010110";
    constant hc_166 : std_logic_vector (7 downto 0) := "00010101";
    signal hc_168 : std_logic_vector (7 downto 0);
    signal hc_172 : std_logic_vector (7 downto 0);
    constant hc_163 : std_logic_vector (7 downto 0) := "00010100";
    constant hc_162 : std_logic_vector (7 downto 0) := "00010011";
    signal hc_164 : std_logic_vector (7 downto 0);
    constant hc_160 : std_logic_vector (7 downto 0) := "00010010";
    constant hc_159 : std_logic_vector (7 downto 0) := "00010001";
    signal hc_161 : std_logic_vector (7 downto 0);
    signal hc_165 : std_logic_vector (7 downto 0);
    signal hc_173 : std_logic_vector (7 downto 0);
    constant hc_155 : std_logic_vector (7 downto 0) := "00010000";
    constant hc_154 : std_logic_vector (7 downto 0) := "00001111";
    signal hc_156 : std_logic_vector (7 downto 0);
    constant hc_152 : std_logic_vector (7 downto 0) := "00001110";
    constant hc_151 : std_logic_vector (7 downto 0) := "00001101";
    signal hc_153 : std_logic_vector (7 downto 0);
    signal hc_157 : std_logic_vector (7 downto 0);
    constant hc_148 : std_logic_vector (7 downto 0) := "00001100";
    constant hc_147 : std_logic_vector (7 downto 0) := "00001011";
    signal hc_149 : std_logic_vector (7 downto 0);
    constant hc_145 : std_logic_vector (7 downto 0) := "00001010";
    constant hc_144 : std_logic_vector (7 downto 0) := "00001001";
    signal hc_146 : std_logic_vector (7 downto 0);
    signal hc_150 : std_logic_vector (7 downto 0);
    signal hc_158 : std_logic_vector (7 downto 0);
    signal hc_174 : std_logic_vector (7 downto 0);
    constant hc_140 : std_logic_vector (7 downto 0) := "00001000";
    constant hc_139 : std_logic_vector (7 downto 0) := "00000111";
    signal hc_141 : std_logic_vector (7 downto 0);
    constant hc_137 : std_logic_vector (7 downto 0) := "00000110";
    constant hc_136 : std_logic_vector (7 downto 0) := "00000101";
    signal hc_138 : std_logic_vector (7 downto 0);
    signal hc_142 : std_logic_vector (7 downto 0);
    constant hc_133 : std_logic_vector (7 downto 0) := "00000100";
    constant hc_132 : std_logic_vector (7 downto 0) := "00000011";
    signal hc_134 : std_logic_vector (7 downto 0);
    constant hc_130 : std_logic_vector (7 downto 0) := "00000010";
    constant hc_129 : std_logic_vector (7 downto 0) := "00000001";
    signal hc_131 : std_logic_vector (7 downto 0);
    signal hc_135 : std_logic_vector (7 downto 0);
    signal hc_143 : std_logic_vector (7 downto 0);
    signal hc_175 : std_logic_vector (7 downto 0);
    constant hc_128 : std_logic_vector (7 downto 0) := "00000000";
    signal hc_123 : std_logic;
    signal hc_122 : std_logic;
    signal hc_124 : std_logic;
    signal hc_120 : std_logic;
    signal hc_119 : std_logic;
    signal hc_121 : std_logic;
    signal hc_125 : std_logic;
    signal hc_116 : std_logic;
    signal hc_115 : std_logic;
    signal hc_117 : std_logic;
    signal hc_113 : std_logic;
    signal hc_112 : std_logic;
    signal hc_114 : std_logic;
    signal hc_118 : std_logic;
    signal hc_126 : std_logic;
    signal hc_107 : std_logic;
    signal hc_106 : std_logic;
    signal hc_108 : std_logic;
    signal hc_104 : std_logic;
    signal hc_103 : std_logic;
    signal hc_105 : std_logic;
    signal hc_109 : std_logic;
    signal hc_100 : std_logic;
    signal hc_99 : std_logic;
    signal hc_101 : std_logic;
    signal hc_97 : std_logic;
    signal hc_96 : std_logic;
    signal hc_98 : std_logic;
    signal hc_102 : std_logic;
    signal hc_110 : std_logic;
    signal hc_92 : std_logic;
    signal hc_91 : std_logic;
    signal hc_93 : std_logic;
    signal hc_89 : std_logic;
    signal hc_88 : std_logic;
    signal hc_90 : std_logic;
    signal hc_94 : std_logic;
    signal hc_85 : std_logic;
    signal hc_84 : std_logic;
    signal hc_86 : std_logic;
    signal hc_82 : std_logic;
    signal hc_79 : std_logic;
    signal hc_78 : std_logic;
    signal hc_77 : std_logic;
    signal hc_76 : std_logic;
    signal hc_75 : std_logic;
    signal hc_74 : std_logic;
    signal hc_73 : std_logic;
    signal hc_72 : std_logic;
    signal hc_71 : std_logic;
    signal hc_70 : std_logic;
    signal hc_69 : std_logic;
    signal hc_68 : std_logic;
    signal hc_67 : std_logic;
    signal hc_66 : std_logic;
    signal hc_65 : std_logic;
    signal hc_64 : std_logic;
    signal hc_63 : std_logic;
    signal hc_62 : std_logic;
    signal hc_61 : std_logic;
    signal hc_60 : std_logic;
    signal hc_59 : std_logic;
    signal hc_58 : std_logic;
    signal hc_57 : std_logic;
    signal hc_52 : std_logic;
    signal hc_53 : std_logic;
    signal hc_50 : std_logic;
    signal hc_51 : std_logic;
    signal hc_48 : std_logic;
    signal hc_49 : std_logic;
    signal hc_46 : std_logic;
    signal hc_47 : std_logic;
    signal hc_44 : std_logic;
    signal hc_45 : std_logic;
    signal hc_42 : std_logic;
    signal hc_43 : std_logic;
    signal hc_40 : std_logic;
    signal hc_41 : std_logic;
    signal hc_38 : std_logic;
    signal hc_39 : std_logic;
    signal hc_36 : std_logic;
    signal hc_37 : std_logic;
    signal hc_34 : std_logic;
    signal hc_35 : std_logic;
    signal hc_32 : std_logic;
    signal hc_33 : std_logic;
    signal hc_30 : std_logic;
    signal hc_31 : std_logic;
    signal hc_28 : std_logic;
    signal hc_29 : std_logic;
    signal hc_26 : std_logic;
    signal hc_27 : std_logic;
    signal hc_24 : std_logic;
    signal hc_25 : std_logic;
    signal hc_22 : std_logic;
    signal hc_23 : std_logic;
    signal hc_20 : std_logic;
    signal hc_21 : std_logic;
    signal hc_18 : std_logic;
    signal hc_19 : std_logic;
    signal hc_16 : std_logic;
    signal hc_17 : std_logic;
    signal hc_14 : std_logic;
    signal hc_15 : std_logic;
    signal hc_12 : std_logic;
    signal hc_13 : std_logic;
    signal hc_10 : std_logic;
    signal hc_11 : std_logic;
    signal hc_8 : std_logic;
    signal hc_9 : std_logic;
    constant hc_4 : std_logic_vector (23 downto 0) := "000000000000000000000001";
    signal hc_5 : std_logic_vector (23 downto 0);
    signal hc_6 : std_logic;
    signal hc_7 : std_logic;
    signal hc_54 : std_logic_vector (23 downto 0);
    signal hc_3 : std_logic;
    signal hc_55 : std_logic_vector (23 downto 0);
    signal hc_56 : std_logic;
    signal hc_80 : std_logic_vector (23 downto 0);
    signal hc_81 : std_logic;
    signal hc_83 : std_logic;
    signal hc_87 : std_logic;
    signal hc_95 : std_logic;
    signal hc_111 : std_logic;
    signal hc_127 : std_logic;
    signal hc_176 : std_logic_vector (7 downto 0);
    signal hc_178 : std_logic;
    signal hc_936 : std_logic_vector (31 downto 0);

begin

    -- logic
    hc_933 <= hc_sl(hc_910(0 downto 0));
    hc_932 <= hc_sl(hc_910(1 downto 1));
    hc_931 <= hc_sl(hc_910(2 downto 2));
    hc_930 <= hc_sl(hc_910(3 downto 3));
    hc_929 <= hc_sl(hc_910(4 downto 4));
    hc_928 <= hc_sl(hc_910(5 downto 5));
    hc_927 <= hc_sl(hc_910(6 downto 6));
    hc_926 <= hc_sl(hc_910(7 downto 7));
    hc_925 <= hc_sl(hc_910(8 downto 8));
    hc_924 <= hc_sl(hc_910(9 downto 9));
    hc_923 <= hc_sl(hc_910(10 downto 10));
    hc_922 <= hc_sl(hc_910(11 downto 11));
    hc_921 <= hc_sl(hc_910(12 downto 12));
    hc_920 <= hc_sl(hc_910(13 downto 13));
    hc_919 <= hc_sl(hc_910(14 downto 14));
    hc_918 <= hc_sl(hc_910(15 downto 15));
    hc_917 <= hc_sl(hc_910(16 downto 16));
    hc_916 <= hc_sl(hc_910(17 downto 17));
    hc_915 <= hc_sl(hc_910(18 downto 18));
    hc_914 <= hc_sl(hc_910(19 downto 19));
    hc_913 <= hc_sl(hc_910(20 downto 20));
    hc_912 <= hc_sl(hc_910(21 downto 21));
    hc_903 <= hc_sl(hc_880(1 downto 1));
    hc_902 <= hc_sl(hc_880(2 downto 2));
    hc_901 <= hc_sl(hc_880(3 downto 3));
    hc_900 <= hc_sl(hc_880(4 downto 4));
    hc_899 <= hc_sl(hc_880(5 downto 5));
    hc_898 <= hc_sl(hc_880(6 downto 6));
    hc_897 <= hc_sl(hc_880(7 downto 7));
    hc_896 <= hc_sl(hc_880(8 downto 8));
    hc_895 <= hc_sl(hc_880(9 downto 9));
    hc_894 <= hc_sl(hc_880(10 downto 10));
    hc_893 <= hc_sl(hc_880(11 downto 11));
    hc_892 <= hc_sl(hc_880(12 downto 12));
    hc_891 <= hc_sl(hc_880(13 downto 13));
    hc_890 <= hc_sl(hc_880(14 downto 14));
    hc_889 <= hc_sl(hc_880(15 downto 15));
    hc_888 <= hc_sl(hc_880(16 downto 16));
    hc_887 <= hc_sl(hc_880(17 downto 17));
    hc_886 <= hc_sl(hc_880(18 downto 18));
    hc_885 <= hc_sl(hc_880(19 downto 19));
    hc_884 <= hc_sl(hc_880(20 downto 20));
    hc_883 <= hc_sl(hc_880(21 downto 21));
    hc_882 <= hc_sl(hc_880(22 downto 22));
    hc_878 <= hc_55(22 downto 0);
    hc_880 <= hc_878 & hc_879;
    hc_881 <= hc_sl(hc_880(23 downto 23));
    hc_904 <= hc_881 & hc_882 & hc_883 & hc_884 & hc_885 & hc_886 & hc_887 & hc_888 & hc_889 & hc_890 & hc_891 & hc_892 & hc_893 & hc_894 & hc_895 & hc_896 & hc_897 & hc_898 & hc_899 & hc_900 & hc_901 & hc_902 & hc_903;
    hc_876 <= hc_sl(hc_853(1 downto 1));
    hc_875 <= hc_sl(hc_853(2 downto 2));
    hc_874 <= hc_sl(hc_853(3 downto 3));
    hc_873 <= hc_sl(hc_853(4 downto 4));
    hc_872 <= hc_sl(hc_853(5 downto 5));
    hc_871 <= hc_sl(hc_853(6 downto 6));
    hc_870 <= hc_sl(hc_853(7 downto 7));
    hc_869 <= hc_sl(hc_853(8 downto 8));
    hc_868 <= hc_sl(hc_853(9 downto 9));
    hc_867 <= hc_sl(hc_853(10 downto 10));
    hc_866 <= hc_sl(hc_853(11 downto 11));
    hc_865 <= hc_sl(hc_853(12 downto 12));
    hc_864 <= hc_sl(hc_853(13 downto 13));
    hc_863 <= hc_sl(hc_853(14 downto 14));
    hc_862 <= hc_sl(hc_853(15 downto 15));
    hc_861 <= hc_sl(hc_853(16 downto 16));
    hc_860 <= hc_sl(hc_853(17 downto 17));
    hc_859 <= hc_sl(hc_853(18 downto 18));
    hc_858 <= hc_sl(hc_853(19 downto 19));
    hc_857 <= hc_sl(hc_853(20 downto 20));
    hc_856 <= hc_sl(hc_853(21 downto 21));
    hc_855 <= hc_sl(hc_853(22 downto 22));
    hc_851 <= hc_55(21 downto 0);
    hc_853 <= hc_851 & hc_852;
    hc_854 <= hc_sl(hc_853(23 downto 23));
    hc_877 <= hc_854 & hc_855 & hc_856 & hc_857 & hc_858 & hc_859 & hc_860 & hc_861 & hc_862 & hc_863 & hc_864 & hc_865 & hc_866 & hc_867 & hc_868 & hc_869 & hc_870 & hc_871 & hc_872 & hc_873 & hc_874 & hc_875 & hc_876;
    with to_integer(hc_uns(hc_217)) select hc_905 <= 
        hc_877 when 0,
        hc_904 when others;
    hc_848 <= hc_sl(hc_825(1 downto 1));
    hc_847 <= hc_sl(hc_825(2 downto 2));
    hc_846 <= hc_sl(hc_825(3 downto 3));
    hc_845 <= hc_sl(hc_825(4 downto 4));
    hc_844 <= hc_sl(hc_825(5 downto 5));
    hc_843 <= hc_sl(hc_825(6 downto 6));
    hc_842 <= hc_sl(hc_825(7 downto 7));
    hc_841 <= hc_sl(hc_825(8 downto 8));
    hc_840 <= hc_sl(hc_825(9 downto 9));
    hc_839 <= hc_sl(hc_825(10 downto 10));
    hc_838 <= hc_sl(hc_825(11 downto 11));
    hc_837 <= hc_sl(hc_825(12 downto 12));
    hc_836 <= hc_sl(hc_825(13 downto 13));
    hc_835 <= hc_sl(hc_825(14 downto 14));
    hc_834 <= hc_sl(hc_825(15 downto 15));
    hc_833 <= hc_sl(hc_825(16 downto 16));
    hc_832 <= hc_sl(hc_825(17 downto 17));
    hc_831 <= hc_sl(hc_825(18 downto 18));
    hc_830 <= hc_sl(hc_825(19 downto 19));
    hc_829 <= hc_sl(hc_825(20 downto 20));
    hc_828 <= hc_sl(hc_825(21 downto 21));
    hc_827 <= hc_sl(hc_825(22 downto 22));
    hc_823 <= hc_55(20 downto 0);
    hc_825 <= hc_823 & hc_824;
    hc_826 <= hc_sl(hc_825(23 downto 23));
    hc_849 <= hc_826 & hc_827 & hc_828 & hc_829 & hc_830 & hc_831 & hc_832 & hc_833 & hc_834 & hc_835 & hc_836 & hc_837 & hc_838 & hc_839 & hc_840 & hc_841 & hc_842 & hc_843 & hc_844 & hc_845 & hc_846 & hc_847 & hc_848;
    hc_821 <= hc_sl(hc_798(1 downto 1));
    hc_820 <= hc_sl(hc_798(2 downto 2));
    hc_819 <= hc_sl(hc_798(3 downto 3));
    hc_818 <= hc_sl(hc_798(4 downto 4));
    hc_817 <= hc_sl(hc_798(5 downto 5));
    hc_816 <= hc_sl(hc_798(6 downto 6));
    hc_815 <= hc_sl(hc_798(7 downto 7));
    hc_814 <= hc_sl(hc_798(8 downto 8));
    hc_813 <= hc_sl(hc_798(9 downto 9));
    hc_812 <= hc_sl(hc_798(10 downto 10));
    hc_811 <= hc_sl(hc_798(11 downto 11));
    hc_810 <= hc_sl(hc_798(12 downto 12));
    hc_809 <= hc_sl(hc_798(13 downto 13));
    hc_808 <= hc_sl(hc_798(14 downto 14));
    hc_807 <= hc_sl(hc_798(15 downto 15));
    hc_806 <= hc_sl(hc_798(16 downto 16));
    hc_805 <= hc_sl(hc_798(17 downto 17));
    hc_804 <= hc_sl(hc_798(18 downto 18));
    hc_803 <= hc_sl(hc_798(19 downto 19));
    hc_802 <= hc_sl(hc_798(20 downto 20));
    hc_801 <= hc_sl(hc_798(21 downto 21));
    hc_800 <= hc_sl(hc_798(22 downto 22));
    hc_796 <= hc_55(19 downto 0);
    hc_798 <= hc_796 & hc_797;
    hc_799 <= hc_sl(hc_798(23 downto 23));
    hc_822 <= hc_799 & hc_800 & hc_801 & hc_802 & hc_803 & hc_804 & hc_805 & hc_806 & hc_807 & hc_808 & hc_809 & hc_810 & hc_811 & hc_812 & hc_813 & hc_814 & hc_815 & hc_816 & hc_817 & hc_818 & hc_819 & hc_820 & hc_821;
    with to_integer(hc_uns(hc_220)) select hc_850 <= 
        hc_822 when 0,
        hc_849 when others;
    with to_integer(hc_uns(hc_219)) select hc_906 <= 
        hc_850 when 0,
        hc_905 when others;
    hc_792 <= hc_sl(hc_769(1 downto 1));
    hc_791 <= hc_sl(hc_769(2 downto 2));
    hc_790 <= hc_sl(hc_769(3 downto 3));
    hc_789 <= hc_sl(hc_769(4 downto 4));
    hc_788 <= hc_sl(hc_769(5 downto 5));
    hc_787 <= hc_sl(hc_769(6 downto 6));
    hc_786 <= hc_sl(hc_769(7 downto 7));
    hc_785 <= hc_sl(hc_769(8 downto 8));
    hc_784 <= hc_sl(hc_769(9 downto 9));
    hc_783 <= hc_sl(hc_769(10 downto 10));
    hc_782 <= hc_sl(hc_769(11 downto 11));
    hc_781 <= hc_sl(hc_769(12 downto 12));
    hc_780 <= hc_sl(hc_769(13 downto 13));
    hc_779 <= hc_sl(hc_769(14 downto 14));
    hc_778 <= hc_sl(hc_769(15 downto 15));
    hc_777 <= hc_sl(hc_769(16 downto 16));
    hc_776 <= hc_sl(hc_769(17 downto 17));
    hc_775 <= hc_sl(hc_769(18 downto 18));
    hc_774 <= hc_sl(hc_769(19 downto 19));
    hc_773 <= hc_sl(hc_769(20 downto 20));
    hc_772 <= hc_sl(hc_769(21 downto 21));
    hc_771 <= hc_sl(hc_769(22 downto 22));
    hc_767 <= hc_55(18 downto 0);
    hc_769 <= hc_767 & hc_768;
    hc_770 <= hc_sl(hc_769(23 downto 23));
    hc_793 <= hc_770 & hc_771 & hc_772 & hc_773 & hc_774 & hc_775 & hc_776 & hc_777 & hc_778 & hc_779 & hc_780 & hc_781 & hc_782 & hc_783 & hc_784 & hc_785 & hc_786 & hc_787 & hc_788 & hc_789 & hc_790 & hc_791 & hc_792;
    hc_765 <= hc_sl(hc_742(1 downto 1));
    hc_764 <= hc_sl(hc_742(2 downto 2));
    hc_763 <= hc_sl(hc_742(3 downto 3));
    hc_762 <= hc_sl(hc_742(4 downto 4));
    hc_761 <= hc_sl(hc_742(5 downto 5));
    hc_760 <= hc_sl(hc_742(6 downto 6));
    hc_759 <= hc_sl(hc_742(7 downto 7));
    hc_758 <= hc_sl(hc_742(8 downto 8));
    hc_757 <= hc_sl(hc_742(9 downto 9));
    hc_756 <= hc_sl(hc_742(10 downto 10));
    hc_755 <= hc_sl(hc_742(11 downto 11));
    hc_754 <= hc_sl(hc_742(12 downto 12));
    hc_753 <= hc_sl(hc_742(13 downto 13));
    hc_752 <= hc_sl(hc_742(14 downto 14));
    hc_751 <= hc_sl(hc_742(15 downto 15));
    hc_750 <= hc_sl(hc_742(16 downto 16));
    hc_749 <= hc_sl(hc_742(17 downto 17));
    hc_748 <= hc_sl(hc_742(18 downto 18));
    hc_747 <= hc_sl(hc_742(19 downto 19));
    hc_746 <= hc_sl(hc_742(20 downto 20));
    hc_745 <= hc_sl(hc_742(21 downto 21));
    hc_744 <= hc_sl(hc_742(22 downto 22));
    hc_740 <= hc_55(17 downto 0);
    hc_742 <= hc_740 & hc_741;
    hc_743 <= hc_sl(hc_742(23 downto 23));
    hc_766 <= hc_743 & hc_744 & hc_745 & hc_746 & hc_747 & hc_748 & hc_749 & hc_750 & hc_751 & hc_752 & hc_753 & hc_754 & hc_755 & hc_756 & hc_757 & hc_758 & hc_759 & hc_760 & hc_761 & hc_762 & hc_763 & hc_764 & hc_765;
    with to_integer(hc_uns(hc_224)) select hc_794 <= 
        hc_766 when 0,
        hc_793 when others;
    hc_737 <= hc_sl(hc_714(1 downto 1));
    hc_736 <= hc_sl(hc_714(2 downto 2));
    hc_735 <= hc_sl(hc_714(3 downto 3));
    hc_734 <= hc_sl(hc_714(4 downto 4));
    hc_733 <= hc_sl(hc_714(5 downto 5));
    hc_732 <= hc_sl(hc_714(6 downto 6));
    hc_731 <= hc_sl(hc_714(7 downto 7));
    hc_730 <= hc_sl(hc_714(8 downto 8));
    hc_729 <= hc_sl(hc_714(9 downto 9));
    hc_728 <= hc_sl(hc_714(10 downto 10));
    hc_727 <= hc_sl(hc_714(11 downto 11));
    hc_726 <= hc_sl(hc_714(12 downto 12));
    hc_725 <= hc_sl(hc_714(13 downto 13));
    hc_724 <= hc_sl(hc_714(14 downto 14));
    hc_723 <= hc_sl(hc_714(15 downto 15));
    hc_722 <= hc_sl(hc_714(16 downto 16));
    hc_721 <= hc_sl(hc_714(17 downto 17));
    hc_720 <= hc_sl(hc_714(18 downto 18));
    hc_719 <= hc_sl(hc_714(19 downto 19));
    hc_718 <= hc_sl(hc_714(20 downto 20));
    hc_717 <= hc_sl(hc_714(21 downto 21));
    hc_716 <= hc_sl(hc_714(22 downto 22));
    hc_712 <= hc_55(16 downto 0);
    hc_714 <= hc_712 & hc_713;
    hc_715 <= hc_sl(hc_714(23 downto 23));
    hc_738 <= hc_715 & hc_716 & hc_717 & hc_718 & hc_719 & hc_720 & hc_721 & hc_722 & hc_723 & hc_724 & hc_725 & hc_726 & hc_727 & hc_728 & hc_729 & hc_730 & hc_731 & hc_732 & hc_733 & hc_734 & hc_735 & hc_736 & hc_737;
    hc_710 <= hc_sl(hc_687(1 downto 1));
    hc_709 <= hc_sl(hc_687(2 downto 2));
    hc_708 <= hc_sl(hc_687(3 downto 3));
    hc_707 <= hc_sl(hc_687(4 downto 4));
    hc_706 <= hc_sl(hc_687(5 downto 5));
    hc_705 <= hc_sl(hc_687(6 downto 6));
    hc_704 <= hc_sl(hc_687(7 downto 7));
    hc_703 <= hc_sl(hc_687(8 downto 8));
    hc_702 <= hc_sl(hc_687(9 downto 9));
    hc_701 <= hc_sl(hc_687(10 downto 10));
    hc_700 <= hc_sl(hc_687(11 downto 11));
    hc_699 <= hc_sl(hc_687(12 downto 12));
    hc_698 <= hc_sl(hc_687(13 downto 13));
    hc_697 <= hc_sl(hc_687(14 downto 14));
    hc_696 <= hc_sl(hc_687(15 downto 15));
    hc_695 <= hc_sl(hc_687(16 downto 16));
    hc_694 <= hc_sl(hc_687(17 downto 17));
    hc_693 <= hc_sl(hc_687(18 downto 18));
    hc_692 <= hc_sl(hc_687(19 downto 19));
    hc_691 <= hc_sl(hc_687(20 downto 20));
    hc_690 <= hc_sl(hc_687(21 downto 21));
    hc_689 <= hc_sl(hc_687(22 downto 22));
    hc_685 <= hc_55(15 downto 0);
    hc_687 <= hc_685 & hc_686;
    hc_688 <= hc_sl(hc_687(23 downto 23));
    hc_711 <= hc_688 & hc_689 & hc_690 & hc_691 & hc_692 & hc_693 & hc_694 & hc_695 & hc_696 & hc_697 & hc_698 & hc_699 & hc_700 & hc_701 & hc_702 & hc_703 & hc_704 & hc_705 & hc_706 & hc_707 & hc_708 & hc_709 & hc_710;
    with to_integer(hc_uns(hc_227)) select hc_739 <= 
        hc_711 when 0,
        hc_738 when others;
    with to_integer(hc_uns(hc_226)) select hc_795 <= 
        hc_739 when 0,
        hc_794 when others;
    with to_integer(hc_uns(hc_223)) select hc_907 <= 
        hc_795 when 0,
        hc_906 when others;
    hc_680 <= hc_sl(hc_657(1 downto 1));
    hc_679 <= hc_sl(hc_657(2 downto 2));
    hc_678 <= hc_sl(hc_657(3 downto 3));
    hc_677 <= hc_sl(hc_657(4 downto 4));
    hc_676 <= hc_sl(hc_657(5 downto 5));
    hc_675 <= hc_sl(hc_657(6 downto 6));
    hc_674 <= hc_sl(hc_657(7 downto 7));
    hc_673 <= hc_sl(hc_657(8 downto 8));
    hc_672 <= hc_sl(hc_657(9 downto 9));
    hc_671 <= hc_sl(hc_657(10 downto 10));
    hc_670 <= hc_sl(hc_657(11 downto 11));
    hc_669 <= hc_sl(hc_657(12 downto 12));
    hc_668 <= hc_sl(hc_657(13 downto 13));
    hc_667 <= hc_sl(hc_657(14 downto 14));
    hc_666 <= hc_sl(hc_657(15 downto 15));
    hc_665 <= hc_sl(hc_657(16 downto 16));
    hc_664 <= hc_sl(hc_657(17 downto 17));
    hc_663 <= hc_sl(hc_657(18 downto 18));
    hc_662 <= hc_sl(hc_657(19 downto 19));
    hc_661 <= hc_sl(hc_657(20 downto 20));
    hc_660 <= hc_sl(hc_657(21 downto 21));
    hc_659 <= hc_sl(hc_657(22 downto 22));
    hc_655 <= hc_55(14 downto 0);
    hc_657 <= hc_655 & hc_656;
    hc_658 <= hc_sl(hc_657(23 downto 23));
    hc_681 <= hc_658 & hc_659 & hc_660 & hc_661 & hc_662 & hc_663 & hc_664 & hc_665 & hc_666 & hc_667 & hc_668 & hc_669 & hc_670 & hc_671 & hc_672 & hc_673 & hc_674 & hc_675 & hc_676 & hc_677 & hc_678 & hc_679 & hc_680;
    hc_653 <= hc_sl(hc_630(1 downto 1));
    hc_652 <= hc_sl(hc_630(2 downto 2));
    hc_651 <= hc_sl(hc_630(3 downto 3));
    hc_650 <= hc_sl(hc_630(4 downto 4));
    hc_649 <= hc_sl(hc_630(5 downto 5));
    hc_648 <= hc_sl(hc_630(6 downto 6));
    hc_647 <= hc_sl(hc_630(7 downto 7));
    hc_646 <= hc_sl(hc_630(8 downto 8));
    hc_645 <= hc_sl(hc_630(9 downto 9));
    hc_644 <= hc_sl(hc_630(10 downto 10));
    hc_643 <= hc_sl(hc_630(11 downto 11));
    hc_642 <= hc_sl(hc_630(12 downto 12));
    hc_641 <= hc_sl(hc_630(13 downto 13));
    hc_640 <= hc_sl(hc_630(14 downto 14));
    hc_639 <= hc_sl(hc_630(15 downto 15));
    hc_638 <= hc_sl(hc_630(16 downto 16));
    hc_637 <= hc_sl(hc_630(17 downto 17));
    hc_636 <= hc_sl(hc_630(18 downto 18));
    hc_635 <= hc_sl(hc_630(19 downto 19));
    hc_634 <= hc_sl(hc_630(20 downto 20));
    hc_633 <= hc_sl(hc_630(21 downto 21));
    hc_632 <= hc_sl(hc_630(22 downto 22));
    hc_628 <= hc_55(13 downto 0);
    hc_630 <= hc_628 & hc_629;
    hc_631 <= hc_sl(hc_630(23 downto 23));
    hc_654 <= hc_631 & hc_632 & hc_633 & hc_634 & hc_635 & hc_636 & hc_637 & hc_638 & hc_639 & hc_640 & hc_641 & hc_642 & hc_643 & hc_644 & hc_645 & hc_646 & hc_647 & hc_648 & hc_649 & hc_650 & hc_651 & hc_652 & hc_653;
    with to_integer(hc_uns(hc_232)) select hc_682 <= 
        hc_654 when 0,
        hc_681 when others;
    hc_625 <= hc_sl(hc_602(1 downto 1));
    hc_624 <= hc_sl(hc_602(2 downto 2));
    hc_623 <= hc_sl(hc_602(3 downto 3));
    hc_622 <= hc_sl(hc_602(4 downto 4));
    hc_621 <= hc_sl(hc_602(5 downto 5));
    hc_620 <= hc_sl(hc_602(6 downto 6));
    hc_619 <= hc_sl(hc_602(7 downto 7));
    hc_618 <= hc_sl(hc_602(8 downto 8));
    hc_617 <= hc_sl(hc_602(9 downto 9));
    hc_616 <= hc_sl(hc_602(10 downto 10));
    hc_615 <= hc_sl(hc_602(11 downto 11));
    hc_614 <= hc_sl(hc_602(12 downto 12));
    hc_613 <= hc_sl(hc_602(13 downto 13));
    hc_612 <= hc_sl(hc_602(14 downto 14));
    hc_611 <= hc_sl(hc_602(15 downto 15));
    hc_610 <= hc_sl(hc_602(16 downto 16));
    hc_609 <= hc_sl(hc_602(17 downto 17));
    hc_608 <= hc_sl(hc_602(18 downto 18));
    hc_607 <= hc_sl(hc_602(19 downto 19));
    hc_606 <= hc_sl(hc_602(20 downto 20));
    hc_605 <= hc_sl(hc_602(21 downto 21));
    hc_604 <= hc_sl(hc_602(22 downto 22));
    hc_600 <= hc_55(12 downto 0);
    hc_602 <= hc_600 & hc_601;
    hc_603 <= hc_sl(hc_602(23 downto 23));
    hc_626 <= hc_603 & hc_604 & hc_605 & hc_606 & hc_607 & hc_608 & hc_609 & hc_610 & hc_611 & hc_612 & hc_613 & hc_614 & hc_615 & hc_616 & hc_617 & hc_618 & hc_619 & hc_620 & hc_621 & hc_622 & hc_623 & hc_624 & hc_625;
    hc_598 <= hc_sl(hc_575(1 downto 1));
    hc_597 <= hc_sl(hc_575(2 downto 2));
    hc_596 <= hc_sl(hc_575(3 downto 3));
    hc_595 <= hc_sl(hc_575(4 downto 4));
    hc_594 <= hc_sl(hc_575(5 downto 5));
    hc_593 <= hc_sl(hc_575(6 downto 6));
    hc_592 <= hc_sl(hc_575(7 downto 7));
    hc_591 <= hc_sl(hc_575(8 downto 8));
    hc_590 <= hc_sl(hc_575(9 downto 9));
    hc_589 <= hc_sl(hc_575(10 downto 10));
    hc_588 <= hc_sl(hc_575(11 downto 11));
    hc_587 <= hc_sl(hc_575(12 downto 12));
    hc_586 <= hc_sl(hc_575(13 downto 13));
    hc_585 <= hc_sl(hc_575(14 downto 14));
    hc_584 <= hc_sl(hc_575(15 downto 15));
    hc_583 <= hc_sl(hc_575(16 downto 16));
    hc_582 <= hc_sl(hc_575(17 downto 17));
    hc_581 <= hc_sl(hc_575(18 downto 18));
    hc_580 <= hc_sl(hc_575(19 downto 19));
    hc_579 <= hc_sl(hc_575(20 downto 20));
    hc_578 <= hc_sl(hc_575(21 downto 21));
    hc_577 <= hc_sl(hc_575(22 downto 22));
    hc_573 <= hc_55(11 downto 0);
    hc_575 <= hc_573 & hc_574;
    hc_576 <= hc_sl(hc_575(23 downto 23));
    hc_599 <= hc_576 & hc_577 & hc_578 & hc_579 & hc_580 & hc_581 & hc_582 & hc_583 & hc_584 & hc_585 & hc_586 & hc_587 & hc_588 & hc_589 & hc_590 & hc_591 & hc_592 & hc_593 & hc_594 & hc_595 & hc_596 & hc_597 & hc_598;
    with to_integer(hc_uns(hc_235)) select hc_627 <= 
        hc_599 when 0,
        hc_626 when others;
    with to_integer(hc_uns(hc_234)) select hc_683 <= 
        hc_627 when 0,
        hc_682 when others;
    hc_569 <= hc_sl(hc_546(1 downto 1));
    hc_568 <= hc_sl(hc_546(2 downto 2));
    hc_567 <= hc_sl(hc_546(3 downto 3));
    hc_566 <= hc_sl(hc_546(4 downto 4));
    hc_565 <= hc_sl(hc_546(5 downto 5));
    hc_564 <= hc_sl(hc_546(6 downto 6));
    hc_563 <= hc_sl(hc_546(7 downto 7));
    hc_562 <= hc_sl(hc_546(8 downto 8));
    hc_561 <= hc_sl(hc_546(9 downto 9));
    hc_560 <= hc_sl(hc_546(10 downto 10));
    hc_559 <= hc_sl(hc_546(11 downto 11));
    hc_558 <= hc_sl(hc_546(12 downto 12));
    hc_557 <= hc_sl(hc_546(13 downto 13));
    hc_556 <= hc_sl(hc_546(14 downto 14));
    hc_555 <= hc_sl(hc_546(15 downto 15));
    hc_554 <= hc_sl(hc_546(16 downto 16));
    hc_553 <= hc_sl(hc_546(17 downto 17));
    hc_552 <= hc_sl(hc_546(18 downto 18));
    hc_551 <= hc_sl(hc_546(19 downto 19));
    hc_550 <= hc_sl(hc_546(20 downto 20));
    hc_549 <= hc_sl(hc_546(21 downto 21));
    hc_548 <= hc_sl(hc_546(22 downto 22));
    hc_544 <= hc_55(10 downto 0);
    hc_546 <= hc_544 & hc_545;
    hc_547 <= hc_sl(hc_546(23 downto 23));
    hc_570 <= hc_547 & hc_548 & hc_549 & hc_550 & hc_551 & hc_552 & hc_553 & hc_554 & hc_555 & hc_556 & hc_557 & hc_558 & hc_559 & hc_560 & hc_561 & hc_562 & hc_563 & hc_564 & hc_565 & hc_566 & hc_567 & hc_568 & hc_569;
    hc_542 <= hc_sl(hc_519(1 downto 1));
    hc_541 <= hc_sl(hc_519(2 downto 2));
    hc_540 <= hc_sl(hc_519(3 downto 3));
    hc_539 <= hc_sl(hc_519(4 downto 4));
    hc_538 <= hc_sl(hc_519(5 downto 5));
    hc_537 <= hc_sl(hc_519(6 downto 6));
    hc_536 <= hc_sl(hc_519(7 downto 7));
    hc_535 <= hc_sl(hc_519(8 downto 8));
    hc_534 <= hc_sl(hc_519(9 downto 9));
    hc_533 <= hc_sl(hc_519(10 downto 10));
    hc_532 <= hc_sl(hc_519(11 downto 11));
    hc_531 <= hc_sl(hc_519(12 downto 12));
    hc_530 <= hc_sl(hc_519(13 downto 13));
    hc_529 <= hc_sl(hc_519(14 downto 14));
    hc_528 <= hc_sl(hc_519(15 downto 15));
    hc_527 <= hc_sl(hc_519(16 downto 16));
    hc_526 <= hc_sl(hc_519(17 downto 17));
    hc_525 <= hc_sl(hc_519(18 downto 18));
    hc_524 <= hc_sl(hc_519(19 downto 19));
    hc_523 <= hc_sl(hc_519(20 downto 20));
    hc_522 <= hc_sl(hc_519(21 downto 21));
    hc_521 <= hc_sl(hc_519(22 downto 22));
    hc_517 <= hc_55(9 downto 0);
    hc_519 <= hc_517 & hc_518;
    hc_520 <= hc_sl(hc_519(23 downto 23));
    hc_543 <= hc_520 & hc_521 & hc_522 & hc_523 & hc_524 & hc_525 & hc_526 & hc_527 & hc_528 & hc_529 & hc_530 & hc_531 & hc_532 & hc_533 & hc_534 & hc_535 & hc_536 & hc_537 & hc_538 & hc_539 & hc_540 & hc_541 & hc_542;
    with to_integer(hc_uns(hc_239)) select hc_571 <= 
        hc_543 when 0,
        hc_570 when others;
    hc_514 <= hc_sl(hc_491(1 downto 1));
    hc_513 <= hc_sl(hc_491(2 downto 2));
    hc_512 <= hc_sl(hc_491(3 downto 3));
    hc_511 <= hc_sl(hc_491(4 downto 4));
    hc_510 <= hc_sl(hc_491(5 downto 5));
    hc_509 <= hc_sl(hc_491(6 downto 6));
    hc_508 <= hc_sl(hc_491(7 downto 7));
    hc_507 <= hc_sl(hc_491(8 downto 8));
    hc_506 <= hc_sl(hc_491(9 downto 9));
    hc_505 <= hc_sl(hc_491(10 downto 10));
    hc_504 <= hc_sl(hc_491(11 downto 11));
    hc_503 <= hc_sl(hc_491(12 downto 12));
    hc_502 <= hc_sl(hc_491(13 downto 13));
    hc_501 <= hc_sl(hc_491(14 downto 14));
    hc_500 <= hc_sl(hc_491(15 downto 15));
    hc_499 <= hc_sl(hc_491(16 downto 16));
    hc_498 <= hc_sl(hc_491(17 downto 17));
    hc_497 <= hc_sl(hc_491(18 downto 18));
    hc_496 <= hc_sl(hc_491(19 downto 19));
    hc_495 <= hc_sl(hc_491(20 downto 20));
    hc_494 <= hc_sl(hc_491(21 downto 21));
    hc_493 <= hc_sl(hc_491(22 downto 22));
    hc_489 <= hc_55(8 downto 0);
    hc_491 <= hc_489 & hc_490;
    hc_492 <= hc_sl(hc_491(23 downto 23));
    hc_515 <= hc_492 & hc_493 & hc_494 & hc_495 & hc_496 & hc_497 & hc_498 & hc_499 & hc_500 & hc_501 & hc_502 & hc_503 & hc_504 & hc_505 & hc_506 & hc_507 & hc_508 & hc_509 & hc_510 & hc_511 & hc_512 & hc_513 & hc_514;
    hc_487 <= hc_sl(hc_464(1 downto 1));
    hc_486 <= hc_sl(hc_464(2 downto 2));
    hc_485 <= hc_sl(hc_464(3 downto 3));
    hc_484 <= hc_sl(hc_464(4 downto 4));
    hc_483 <= hc_sl(hc_464(5 downto 5));
    hc_482 <= hc_sl(hc_464(6 downto 6));
    hc_481 <= hc_sl(hc_464(7 downto 7));
    hc_480 <= hc_sl(hc_464(8 downto 8));
    hc_479 <= hc_sl(hc_464(9 downto 9));
    hc_478 <= hc_sl(hc_464(10 downto 10));
    hc_477 <= hc_sl(hc_464(11 downto 11));
    hc_476 <= hc_sl(hc_464(12 downto 12));
    hc_475 <= hc_sl(hc_464(13 downto 13));
    hc_474 <= hc_sl(hc_464(14 downto 14));
    hc_473 <= hc_sl(hc_464(15 downto 15));
    hc_472 <= hc_sl(hc_464(16 downto 16));
    hc_471 <= hc_sl(hc_464(17 downto 17));
    hc_470 <= hc_sl(hc_464(18 downto 18));
    hc_469 <= hc_sl(hc_464(19 downto 19));
    hc_468 <= hc_sl(hc_464(20 downto 20));
    hc_467 <= hc_sl(hc_464(21 downto 21));
    hc_466 <= hc_sl(hc_464(22 downto 22));
    hc_462 <= hc_55(7 downto 0);
    hc_464 <= hc_462 & hc_463;
    hc_465 <= hc_sl(hc_464(23 downto 23));
    hc_488 <= hc_465 & hc_466 & hc_467 & hc_468 & hc_469 & hc_470 & hc_471 & hc_472 & hc_473 & hc_474 & hc_475 & hc_476 & hc_477 & hc_478 & hc_479 & hc_480 & hc_481 & hc_482 & hc_483 & hc_484 & hc_485 & hc_486 & hc_487;
    with to_integer(hc_uns(hc_242)) select hc_516 <= 
        hc_488 when 0,
        hc_515 when others;
    with to_integer(hc_uns(hc_241)) select hc_572 <= 
        hc_516 when 0,
        hc_571 when others;
    with to_integer(hc_uns(hc_238)) select hc_684 <= 
        hc_572 when 0,
        hc_683 when others;
    with to_integer(hc_uns(hc_231)) select hc_908 <= 
        hc_684 when 0,
        hc_907 when others;
    hc_457 <= hc_sl(hc_434(1 downto 1));
    hc_456 <= hc_sl(hc_434(2 downto 2));
    hc_455 <= hc_sl(hc_434(3 downto 3));
    hc_454 <= hc_sl(hc_434(4 downto 4));
    hc_453 <= hc_sl(hc_434(5 downto 5));
    hc_452 <= hc_sl(hc_434(6 downto 6));
    hc_451 <= hc_sl(hc_434(7 downto 7));
    hc_450 <= hc_sl(hc_434(8 downto 8));
    hc_449 <= hc_sl(hc_434(9 downto 9));
    hc_448 <= hc_sl(hc_434(10 downto 10));
    hc_447 <= hc_sl(hc_434(11 downto 11));
    hc_446 <= hc_sl(hc_434(12 downto 12));
    hc_445 <= hc_sl(hc_434(13 downto 13));
    hc_444 <= hc_sl(hc_434(14 downto 14));
    hc_443 <= hc_sl(hc_434(15 downto 15));
    hc_442 <= hc_sl(hc_434(16 downto 16));
    hc_441 <= hc_sl(hc_434(17 downto 17));
    hc_440 <= hc_sl(hc_434(18 downto 18));
    hc_439 <= hc_sl(hc_434(19 downto 19));
    hc_438 <= hc_sl(hc_434(20 downto 20));
    hc_437 <= hc_sl(hc_434(21 downto 21));
    hc_436 <= hc_sl(hc_434(22 downto 22));
    hc_432 <= hc_55(6 downto 0);
    hc_434 <= hc_432 & hc_433;
    hc_435 <= hc_sl(hc_434(23 downto 23));
    hc_458 <= hc_435 & hc_436 & hc_437 & hc_438 & hc_439 & hc_440 & hc_441 & hc_442 & hc_443 & hc_444 & hc_445 & hc_446 & hc_447 & hc_448 & hc_449 & hc_450 & hc_451 & hc_452 & hc_453 & hc_454 & hc_455 & hc_456 & hc_457;
    hc_430 <= hc_sl(hc_407(1 downto 1));
    hc_429 <= hc_sl(hc_407(2 downto 2));
    hc_428 <= hc_sl(hc_407(3 downto 3));
    hc_427 <= hc_sl(hc_407(4 downto 4));
    hc_426 <= hc_sl(hc_407(5 downto 5));
    hc_425 <= hc_sl(hc_407(6 downto 6));
    hc_424 <= hc_sl(hc_407(7 downto 7));
    hc_423 <= hc_sl(hc_407(8 downto 8));
    hc_422 <= hc_sl(hc_407(9 downto 9));
    hc_421 <= hc_sl(hc_407(10 downto 10));
    hc_420 <= hc_sl(hc_407(11 downto 11));
    hc_419 <= hc_sl(hc_407(12 downto 12));
    hc_418 <= hc_sl(hc_407(13 downto 13));
    hc_417 <= hc_sl(hc_407(14 downto 14));
    hc_416 <= hc_sl(hc_407(15 downto 15));
    hc_415 <= hc_sl(hc_407(16 downto 16));
    hc_414 <= hc_sl(hc_407(17 downto 17));
    hc_413 <= hc_sl(hc_407(18 downto 18));
    hc_412 <= hc_sl(hc_407(19 downto 19));
    hc_411 <= hc_sl(hc_407(20 downto 20));
    hc_410 <= hc_sl(hc_407(21 downto 21));
    hc_409 <= hc_sl(hc_407(22 downto 22));
    hc_405 <= hc_55(5 downto 0);
    hc_407 <= hc_405 & hc_406;
    hc_408 <= hc_sl(hc_407(23 downto 23));
    hc_431 <= hc_408 & hc_409 & hc_410 & hc_411 & hc_412 & hc_413 & hc_414 & hc_415 & hc_416 & hc_417 & hc_418 & hc_419 & hc_420 & hc_421 & hc_422 & hc_423 & hc_424 & hc_425 & hc_426 & hc_427 & hc_428 & hc_429 & hc_430;
    with to_integer(hc_uns(hc_248)) select hc_459 <= 
        hc_431 when 0,
        hc_458 when others;
    hc_402 <= hc_sl(hc_379(1 downto 1));
    hc_401 <= hc_sl(hc_379(2 downto 2));
    hc_400 <= hc_sl(hc_379(3 downto 3));
    hc_399 <= hc_sl(hc_379(4 downto 4));
    hc_398 <= hc_sl(hc_379(5 downto 5));
    hc_397 <= hc_sl(hc_379(6 downto 6));
    hc_396 <= hc_sl(hc_379(7 downto 7));
    hc_395 <= hc_sl(hc_379(8 downto 8));
    hc_394 <= hc_sl(hc_379(9 downto 9));
    hc_393 <= hc_sl(hc_379(10 downto 10));
    hc_392 <= hc_sl(hc_379(11 downto 11));
    hc_391 <= hc_sl(hc_379(12 downto 12));
    hc_390 <= hc_sl(hc_379(13 downto 13));
    hc_389 <= hc_sl(hc_379(14 downto 14));
    hc_388 <= hc_sl(hc_379(15 downto 15));
    hc_387 <= hc_sl(hc_379(16 downto 16));
    hc_386 <= hc_sl(hc_379(17 downto 17));
    hc_385 <= hc_sl(hc_379(18 downto 18));
    hc_384 <= hc_sl(hc_379(19 downto 19));
    hc_383 <= hc_sl(hc_379(20 downto 20));
    hc_382 <= hc_sl(hc_379(21 downto 21));
    hc_381 <= hc_sl(hc_379(22 downto 22));
    hc_377 <= hc_55(4 downto 0);
    hc_379 <= hc_377 & hc_378;
    hc_380 <= hc_sl(hc_379(23 downto 23));
    hc_403 <= hc_380 & hc_381 & hc_382 & hc_383 & hc_384 & hc_385 & hc_386 & hc_387 & hc_388 & hc_389 & hc_390 & hc_391 & hc_392 & hc_393 & hc_394 & hc_395 & hc_396 & hc_397 & hc_398 & hc_399 & hc_400 & hc_401 & hc_402;
    hc_375 <= hc_sl(hc_352(1 downto 1));
    hc_374 <= hc_sl(hc_352(2 downto 2));
    hc_373 <= hc_sl(hc_352(3 downto 3));
    hc_372 <= hc_sl(hc_352(4 downto 4));
    hc_371 <= hc_sl(hc_352(5 downto 5));
    hc_370 <= hc_sl(hc_352(6 downto 6));
    hc_369 <= hc_sl(hc_352(7 downto 7));
    hc_368 <= hc_sl(hc_352(8 downto 8));
    hc_367 <= hc_sl(hc_352(9 downto 9));
    hc_366 <= hc_sl(hc_352(10 downto 10));
    hc_365 <= hc_sl(hc_352(11 downto 11));
    hc_364 <= hc_sl(hc_352(12 downto 12));
    hc_363 <= hc_sl(hc_352(13 downto 13));
    hc_362 <= hc_sl(hc_352(14 downto 14));
    hc_361 <= hc_sl(hc_352(15 downto 15));
    hc_360 <= hc_sl(hc_352(16 downto 16));
    hc_359 <= hc_sl(hc_352(17 downto 17));
    hc_358 <= hc_sl(hc_352(18 downto 18));
    hc_357 <= hc_sl(hc_352(19 downto 19));
    hc_356 <= hc_sl(hc_352(20 downto 20));
    hc_355 <= hc_sl(hc_352(21 downto 21));
    hc_354 <= hc_sl(hc_352(22 downto 22));
    hc_350 <= hc_55(3 downto 0);
    hc_352 <= hc_350 & hc_351;
    hc_353 <= hc_sl(hc_352(23 downto 23));
    hc_376 <= hc_353 & hc_354 & hc_355 & hc_356 & hc_357 & hc_358 & hc_359 & hc_360 & hc_361 & hc_362 & hc_363 & hc_364 & hc_365 & hc_366 & hc_367 & hc_368 & hc_369 & hc_370 & hc_371 & hc_372 & hc_373 & hc_374 & hc_375;
    with to_integer(hc_uns(hc_251)) select hc_404 <= 
        hc_376 when 0,
        hc_403 when others;
    with to_integer(hc_uns(hc_250)) select hc_460 <= 
        hc_404 when 0,
        hc_459 when others;
    hc_346 <= hc_sl(hc_323(1 downto 1));
    hc_345 <= hc_sl(hc_323(2 downto 2));
    hc_344 <= hc_sl(hc_323(3 downto 3));
    hc_343 <= hc_sl(hc_323(4 downto 4));
    hc_342 <= hc_sl(hc_323(5 downto 5));
    hc_341 <= hc_sl(hc_323(6 downto 6));
    hc_340 <= hc_sl(hc_323(7 downto 7));
    hc_339 <= hc_sl(hc_323(8 downto 8));
    hc_338 <= hc_sl(hc_323(9 downto 9));
    hc_337 <= hc_sl(hc_323(10 downto 10));
    hc_336 <= hc_sl(hc_323(11 downto 11));
    hc_335 <= hc_sl(hc_323(12 downto 12));
    hc_334 <= hc_sl(hc_323(13 downto 13));
    hc_333 <= hc_sl(hc_323(14 downto 14));
    hc_332 <= hc_sl(hc_323(15 downto 15));
    hc_331 <= hc_sl(hc_323(16 downto 16));
    hc_330 <= hc_sl(hc_323(17 downto 17));
    hc_329 <= hc_sl(hc_323(18 downto 18));
    hc_328 <= hc_sl(hc_323(19 downto 19));
    hc_327 <= hc_sl(hc_323(20 downto 20));
    hc_326 <= hc_sl(hc_323(21 downto 21));
    hc_325 <= hc_sl(hc_323(22 downto 22));
    hc_321 <= hc_55(2 downto 0);
    hc_323 <= hc_321 & hc_322;
    hc_324 <= hc_sl(hc_323(23 downto 23));
    hc_347 <= hc_324 & hc_325 & hc_326 & hc_327 & hc_328 & hc_329 & hc_330 & hc_331 & hc_332 & hc_333 & hc_334 & hc_335 & hc_336 & hc_337 & hc_338 & hc_339 & hc_340 & hc_341 & hc_342 & hc_343 & hc_344 & hc_345 & hc_346;
    hc_319 <= hc_sl(hc_296(1 downto 1));
    hc_318 <= hc_sl(hc_296(2 downto 2));
    hc_317 <= hc_sl(hc_296(3 downto 3));
    hc_316 <= hc_sl(hc_296(4 downto 4));
    hc_315 <= hc_sl(hc_296(5 downto 5));
    hc_314 <= hc_sl(hc_296(6 downto 6));
    hc_313 <= hc_sl(hc_296(7 downto 7));
    hc_312 <= hc_sl(hc_296(8 downto 8));
    hc_311 <= hc_sl(hc_296(9 downto 9));
    hc_310 <= hc_sl(hc_296(10 downto 10));
    hc_309 <= hc_sl(hc_296(11 downto 11));
    hc_308 <= hc_sl(hc_296(12 downto 12));
    hc_307 <= hc_sl(hc_296(13 downto 13));
    hc_306 <= hc_sl(hc_296(14 downto 14));
    hc_305 <= hc_sl(hc_296(15 downto 15));
    hc_304 <= hc_sl(hc_296(16 downto 16));
    hc_303 <= hc_sl(hc_296(17 downto 17));
    hc_302 <= hc_sl(hc_296(18 downto 18));
    hc_301 <= hc_sl(hc_296(19 downto 19));
    hc_300 <= hc_sl(hc_296(20 downto 20));
    hc_299 <= hc_sl(hc_296(21 downto 21));
    hc_298 <= hc_sl(hc_296(22 downto 22));
    hc_294 <= hc_55(1 downto 0);
    hc_296 <= hc_294 & hc_295;
    hc_297 <= hc_sl(hc_296(23 downto 23));
    hc_320 <= hc_297 & hc_298 & hc_299 & hc_300 & hc_301 & hc_302 & hc_303 & hc_304 & hc_305 & hc_306 & hc_307 & hc_308 & hc_309 & hc_310 & hc_311 & hc_312 & hc_313 & hc_314 & hc_315 & hc_316 & hc_317 & hc_318 & hc_319;
    with to_integer(hc_uns(hc_255)) select hc_348 <= 
        hc_320 when 0,
        hc_347 when others;
    hc_291 <= hc_sl(hc_268(1 downto 1));
    hc_290 <= hc_sl(hc_268(2 downto 2));
    hc_289 <= hc_sl(hc_268(3 downto 3));
    hc_288 <= hc_sl(hc_268(4 downto 4));
    hc_287 <= hc_sl(hc_268(5 downto 5));
    hc_286 <= hc_sl(hc_268(6 downto 6));
    hc_285 <= hc_sl(hc_268(7 downto 7));
    hc_284 <= hc_sl(hc_268(8 downto 8));
    hc_283 <= hc_sl(hc_268(9 downto 9));
    hc_282 <= hc_sl(hc_268(10 downto 10));
    hc_281 <= hc_sl(hc_268(11 downto 11));
    hc_280 <= hc_sl(hc_268(12 downto 12));
    hc_279 <= hc_sl(hc_268(13 downto 13));
    hc_278 <= hc_sl(hc_268(14 downto 14));
    hc_277 <= hc_sl(hc_268(15 downto 15));
    hc_276 <= hc_sl(hc_268(16 downto 16));
    hc_275 <= hc_sl(hc_268(17 downto 17));
    hc_274 <= hc_sl(hc_268(18 downto 18));
    hc_273 <= hc_sl(hc_268(19 downto 19));
    hc_272 <= hc_sl(hc_268(20 downto 20));
    hc_271 <= hc_sl(hc_268(21 downto 21));
    hc_270 <= hc_sl(hc_268(22 downto 22));
    hc_266 <= hc_sl(hc_55(0 downto 0));
    hc_268 <= hc_266 & hc_267;
    hc_269 <= hc_sl(hc_268(23 downto 23));
    hc_292 <= hc_269 & hc_270 & hc_271 & hc_272 & hc_273 & hc_274 & hc_275 & hc_276 & hc_277 & hc_278 & hc_279 & hc_280 & hc_281 & hc_282 & hc_283 & hc_284 & hc_285 & hc_286 & hc_287 & hc_288 & hc_289 & hc_290 & hc_291;
    with to_integer(hc_uns(hc_258)) select hc_293 <= 
        hc_265 when 0,
        hc_292 when others;
    with to_integer(hc_uns(hc_257)) select hc_349 <= 
        hc_293 when 0,
        hc_348 when others;
    with to_integer(hc_uns(hc_254)) select hc_461 <= 
        hc_349 when 0,
        hc_460 when others;
    with to_integer(hc_uns(hc_247)) select hc_909 <= 
        hc_461 when 0,
        hc_908 when others;
    hc_259 <= hc_sl(hc_216(23 downto 23));
    hc_258 <= hc_sl(hc_216(22 downto 22));
    hc_260 <= hc_sl(hc_uns(hc_258) or hc_uns(hc_259));
    hc_256 <= hc_sl(hc_216(21 downto 21));
    hc_255 <= hc_sl(hc_216(20 downto 20));
    hc_257 <= hc_sl(hc_uns(hc_255) or hc_uns(hc_256));
    hc_261 <= hc_sl(hc_uns(hc_257) or hc_uns(hc_260));
    hc_252 <= hc_sl(hc_216(19 downto 19));
    hc_251 <= hc_sl(hc_216(18 downto 18));
    hc_253 <= hc_sl(hc_uns(hc_251) or hc_uns(hc_252));
    hc_249 <= hc_sl(hc_216(17 downto 17));
    hc_248 <= hc_sl(hc_216(16 downto 16));
    hc_250 <= hc_sl(hc_uns(hc_248) or hc_uns(hc_249));
    hc_254 <= hc_sl(hc_uns(hc_250) or hc_uns(hc_253));
    hc_262 <= hc_sl(hc_uns(hc_254) or hc_uns(hc_261));
    hc_243 <= hc_sl(hc_216(15 downto 15));
    hc_242 <= hc_sl(hc_216(14 downto 14));
    hc_244 <= hc_sl(hc_uns(hc_242) or hc_uns(hc_243));
    hc_240 <= hc_sl(hc_216(13 downto 13));
    hc_239 <= hc_sl(hc_216(12 downto 12));
    hc_241 <= hc_sl(hc_uns(hc_239) or hc_uns(hc_240));
    hc_245 <= hc_sl(hc_uns(hc_241) or hc_uns(hc_244));
    hc_236 <= hc_sl(hc_216(11 downto 11));
    hc_235 <= hc_sl(hc_216(10 downto 10));
    hc_237 <= hc_sl(hc_uns(hc_235) or hc_uns(hc_236));
    hc_233 <= hc_sl(hc_216(9 downto 9));
    hc_232 <= hc_sl(hc_216(8 downto 8));
    hc_234 <= hc_sl(hc_uns(hc_232) or hc_uns(hc_233));
    hc_238 <= hc_sl(hc_uns(hc_234) or hc_uns(hc_237));
    hc_246 <= hc_sl(hc_uns(hc_238) or hc_uns(hc_245));
    hc_228 <= hc_sl(hc_216(7 downto 7));
    hc_227 <= hc_sl(hc_216(6 downto 6));
    hc_229 <= hc_sl(hc_uns(hc_227) or hc_uns(hc_228));
    hc_225 <= hc_sl(hc_216(5 downto 5));
    hc_224 <= hc_sl(hc_216(4 downto 4));
    hc_226 <= hc_sl(hc_uns(hc_224) or hc_uns(hc_225));
    hc_230 <= hc_sl(hc_uns(hc_226) or hc_uns(hc_229));
    hc_221 <= hc_sl(hc_216(3 downto 3));
    hc_220 <= hc_sl(hc_216(2 downto 2));
    hc_222 <= hc_sl(hc_uns(hc_220) or hc_uns(hc_221));
    hc_218 <= hc_sl(hc_216(1 downto 1));
    hc_215 <= hc_sl(hc_55(23 downto 23));
    hc_214 <= hc_sl(hc_55(22 downto 22));
    hc_213 <= hc_sl(hc_55(21 downto 21));
    hc_212 <= hc_sl(hc_55(20 downto 20));
    hc_211 <= hc_sl(hc_55(19 downto 19));
    hc_210 <= hc_sl(hc_55(18 downto 18));
    hc_209 <= hc_sl(hc_55(17 downto 17));
    hc_208 <= hc_sl(hc_55(16 downto 16));
    hc_207 <= hc_sl(hc_55(15 downto 15));
    hc_206 <= hc_sl(hc_55(14 downto 14));
    hc_205 <= hc_sl(hc_55(13 downto 13));
    hc_204 <= hc_sl(hc_55(12 downto 12));
    hc_203 <= hc_sl(hc_55(11 downto 11));
    hc_202 <= hc_sl(hc_55(10 downto 10));
    hc_201 <= hc_sl(hc_55(9 downto 9));
    hc_200 <= hc_sl(hc_55(8 downto 8));
    hc_199 <= hc_sl(hc_55(7 downto 7));
    hc_198 <= hc_sl(hc_55(6 downto 6));
    hc_197 <= hc_sl(hc_55(5 downto 5));
    hc_196 <= hc_sl(hc_55(4 downto 4));
    hc_195 <= hc_sl(hc_55(3 downto 3));
    hc_194 <= hc_sl(hc_55(2 downto 2));
    hc_193 <= hc_sl(hc_55(1 downto 1));
    hc_192 <= hc_sl(hc_55(0 downto 0));
    hc_216 <= hc_192 & hc_193 & hc_194 & hc_195 & hc_196 & hc_197 & hc_198 & hc_199 & hc_200 & hc_201 & hc_202 & hc_203 & hc_204 & hc_205 & hc_206 & hc_207 & hc_208 & hc_209 & hc_210 & hc_211 & hc_212 & hc_213 & hc_214 & hc_215;
    hc_217 <= hc_sl(hc_216(0 downto 0));
    hc_219 <= hc_sl(hc_uns(hc_217) or hc_uns(hc_218));
    hc_223 <= hc_sl(hc_uns(hc_219) or hc_uns(hc_222));
    hc_231 <= hc_sl(hc_uns(hc_223) or hc_uns(hc_230));
    hc_247 <= hc_sl(hc_uns(hc_231) or hc_uns(hc_246));
    hc_263 <= hc_sl(hc_uns(hc_247) or hc_uns(hc_262));
    with to_integer(hc_uns(hc_263)) select hc_910 <= 
        hc_264 when 0,
        hc_909 when others;
    hc_911 <= hc_sl(hc_910(22 downto 22));
    hc_191 <= hc_sl(hc_183(0 downto 0));
    hc_190 <= hc_sl(hc_183(1 downto 1));
    hc_189 <= hc_sl(hc_183(2 downto 2));
    hc_188 <= hc_sl(hc_183(3 downto 3));
    hc_187 <= hc_sl(hc_183(4 downto 4));
    hc_186 <= hc_sl(hc_183(5 downto 5));
    hc_185 <= hc_sl(hc_183(6 downto 6));
    hc_181 <= hc_slv(hc_uns(hc_176) - hc_uns(hc_180));
    hc_183 <= hc_slv(hc_uns(hc_181) + hc_uns(hc_182));
    hc_184 <= hc_sl(hc_183(7 downto 7));
    hc_179 <= hc_sl(a(23 downto 23));
    hc_934 <= hc_179 & hc_184 & hc_185 & hc_186 & hc_187 & hc_188 & hc_189 & hc_190 & hc_191 & hc_911 & hc_912 & hc_913 & hc_914 & hc_915 & hc_916 & hc_917 & hc_918 & hc_919 & hc_920 & hc_921 & hc_922 & hc_923 & hc_924 & hc_925 & hc_926 & hc_927 & hc_928 & hc_929 & hc_930 & hc_931 & hc_932 & hc_933;
    with to_integer(hc_uns(hc_81)) select hc_171 <= 
        hc_169 when 0,
        hc_170 when others;
    with to_integer(hc_uns(hc_84)) select hc_168 <= 
        hc_166 when 0,
        hc_167 when others;
    with to_integer(hc_uns(hc_83)) select hc_172 <= 
        hc_168 when 0,
        hc_171 when others;
    with to_integer(hc_uns(hc_88)) select hc_164 <= 
        hc_162 when 0,
        hc_163 when others;
    with to_integer(hc_uns(hc_91)) select hc_161 <= 
        hc_159 when 0,
        hc_160 when others;
    with to_integer(hc_uns(hc_90)) select hc_165 <= 
        hc_161 when 0,
        hc_164 when others;
    with to_integer(hc_uns(hc_87)) select hc_173 <= 
        hc_165 when 0,
        hc_172 when others;
    with to_integer(hc_uns(hc_96)) select hc_156 <= 
        hc_154 when 0,
        hc_155 when others;
    with to_integer(hc_uns(hc_99)) select hc_153 <= 
        hc_151 when 0,
        hc_152 when others;
    with to_integer(hc_uns(hc_98)) select hc_157 <= 
        hc_153 when 0,
        hc_156 when others;
    with to_integer(hc_uns(hc_103)) select hc_149 <= 
        hc_147 when 0,
        hc_148 when others;
    with to_integer(hc_uns(hc_106)) select hc_146 <= 
        hc_144 when 0,
        hc_145 when others;
    with to_integer(hc_uns(hc_105)) select hc_150 <= 
        hc_146 when 0,
        hc_149 when others;
    with to_integer(hc_uns(hc_102)) select hc_158 <= 
        hc_150 when 0,
        hc_157 when others;
    with to_integer(hc_uns(hc_95)) select hc_174 <= 
        hc_158 when 0,
        hc_173 when others;
    with to_integer(hc_uns(hc_112)) select hc_141 <= 
        hc_139 when 0,
        hc_140 when others;
    with to_integer(hc_uns(hc_115)) select hc_138 <= 
        hc_136 when 0,
        hc_137 when others;
    with to_integer(hc_uns(hc_114)) select hc_142 <= 
        hc_138 when 0,
        hc_141 when others;
    with to_integer(hc_uns(hc_119)) select hc_134 <= 
        hc_132 when 0,
        hc_133 when others;
    with to_integer(hc_uns(hc_122)) select hc_131 <= 
        hc_129 when 0,
        hc_130 when others;
    with to_integer(hc_uns(hc_121)) select hc_135 <= 
        hc_131 when 0,
        hc_134 when others;
    with to_integer(hc_uns(hc_118)) select hc_143 <= 
        hc_135 when 0,
        hc_142 when others;
    with to_integer(hc_uns(hc_111)) select hc_175 <= 
        hc_143 when 0,
        hc_174 when others;
    hc_123 <= hc_sl(hc_80(23 downto 23));
    hc_122 <= hc_sl(hc_80(22 downto 22));
    hc_124 <= hc_sl(hc_uns(hc_122) or hc_uns(hc_123));
    hc_120 <= hc_sl(hc_80(21 downto 21));
    hc_119 <= hc_sl(hc_80(20 downto 20));
    hc_121 <= hc_sl(hc_uns(hc_119) or hc_uns(hc_120));
    hc_125 <= hc_sl(hc_uns(hc_121) or hc_uns(hc_124));
    hc_116 <= hc_sl(hc_80(19 downto 19));
    hc_115 <= hc_sl(hc_80(18 downto 18));
    hc_117 <= hc_sl(hc_uns(hc_115) or hc_uns(hc_116));
    hc_113 <= hc_sl(hc_80(17 downto 17));
    hc_112 <= hc_sl(hc_80(16 downto 16));
    hc_114 <= hc_sl(hc_uns(hc_112) or hc_uns(hc_113));
    hc_118 <= hc_sl(hc_uns(hc_114) or hc_uns(hc_117));
    hc_126 <= hc_sl(hc_uns(hc_118) or hc_uns(hc_125));
    hc_107 <= hc_sl(hc_80(15 downto 15));
    hc_106 <= hc_sl(hc_80(14 downto 14));
    hc_108 <= hc_sl(hc_uns(hc_106) or hc_uns(hc_107));
    hc_104 <= hc_sl(hc_80(13 downto 13));
    hc_103 <= hc_sl(hc_80(12 downto 12));
    hc_105 <= hc_sl(hc_uns(hc_103) or hc_uns(hc_104));
    hc_109 <= hc_sl(hc_uns(hc_105) or hc_uns(hc_108));
    hc_100 <= hc_sl(hc_80(11 downto 11));
    hc_99 <= hc_sl(hc_80(10 downto 10));
    hc_101 <= hc_sl(hc_uns(hc_99) or hc_uns(hc_100));
    hc_97 <= hc_sl(hc_80(9 downto 9));
    hc_96 <= hc_sl(hc_80(8 downto 8));
    hc_98 <= hc_sl(hc_uns(hc_96) or hc_uns(hc_97));
    hc_102 <= hc_sl(hc_uns(hc_98) or hc_uns(hc_101));
    hc_110 <= hc_sl(hc_uns(hc_102) or hc_uns(hc_109));
    hc_92 <= hc_sl(hc_80(7 downto 7));
    hc_91 <= hc_sl(hc_80(6 downto 6));
    hc_93 <= hc_sl(hc_uns(hc_91) or hc_uns(hc_92));
    hc_89 <= hc_sl(hc_80(5 downto 5));
    hc_88 <= hc_sl(hc_80(4 downto 4));
    hc_90 <= hc_sl(hc_uns(hc_88) or hc_uns(hc_89));
    hc_94 <= hc_sl(hc_uns(hc_90) or hc_uns(hc_93));
    hc_85 <= hc_sl(hc_80(3 downto 3));
    hc_84 <= hc_sl(hc_80(2 downto 2));
    hc_86 <= hc_sl(hc_uns(hc_84) or hc_uns(hc_85));
    hc_82 <= hc_sl(hc_80(1 downto 1));
    hc_79 <= hc_sl(hc_55(23 downto 23));
    hc_78 <= hc_sl(hc_55(22 downto 22));
    hc_77 <= hc_sl(hc_55(21 downto 21));
    hc_76 <= hc_sl(hc_55(20 downto 20));
    hc_75 <= hc_sl(hc_55(19 downto 19));
    hc_74 <= hc_sl(hc_55(18 downto 18));
    hc_73 <= hc_sl(hc_55(17 downto 17));
    hc_72 <= hc_sl(hc_55(16 downto 16));
    hc_71 <= hc_sl(hc_55(15 downto 15));
    hc_70 <= hc_sl(hc_55(14 downto 14));
    hc_69 <= hc_sl(hc_55(13 downto 13));
    hc_68 <= hc_sl(hc_55(12 downto 12));
    hc_67 <= hc_sl(hc_55(11 downto 11));
    hc_66 <= hc_sl(hc_55(10 downto 10));
    hc_65 <= hc_sl(hc_55(9 downto 9));
    hc_64 <= hc_sl(hc_55(8 downto 8));
    hc_63 <= hc_sl(hc_55(7 downto 7));
    hc_62 <= hc_sl(hc_55(6 downto 6));
    hc_61 <= hc_sl(hc_55(5 downto 5));
    hc_60 <= hc_sl(hc_55(4 downto 4));
    hc_59 <= hc_sl(hc_55(3 downto 3));
    hc_58 <= hc_sl(hc_55(2 downto 2));
    hc_57 <= hc_sl(hc_55(1 downto 1));
    hc_52 <= hc_sl(hc_5(0 downto 0));
    hc_53 <= hc_sl(not hc_uns(hc_52));
    hc_50 <= hc_sl(hc_5(1 downto 1));
    hc_51 <= hc_sl(not hc_uns(hc_50));
    hc_48 <= hc_sl(hc_5(2 downto 2));
    hc_49 <= hc_sl(not hc_uns(hc_48));
    hc_46 <= hc_sl(hc_5(3 downto 3));
    hc_47 <= hc_sl(not hc_uns(hc_46));
    hc_44 <= hc_sl(hc_5(4 downto 4));
    hc_45 <= hc_sl(not hc_uns(hc_44));
    hc_42 <= hc_sl(hc_5(5 downto 5));
    hc_43 <= hc_sl(not hc_uns(hc_42));
    hc_40 <= hc_sl(hc_5(6 downto 6));
    hc_41 <= hc_sl(not hc_uns(hc_40));
    hc_38 <= hc_sl(hc_5(7 downto 7));
    hc_39 <= hc_sl(not hc_uns(hc_38));
    hc_36 <= hc_sl(hc_5(8 downto 8));
    hc_37 <= hc_sl(not hc_uns(hc_36));
    hc_34 <= hc_sl(hc_5(9 downto 9));
    hc_35 <= hc_sl(not hc_uns(hc_34));
    hc_32 <= hc_sl(hc_5(10 downto 10));
    hc_33 <= hc_sl(not hc_uns(hc_32));
    hc_30 <= hc_sl(hc_5(11 downto 11));
    hc_31 <= hc_sl(not hc_uns(hc_30));
    hc_28 <= hc_sl(hc_5(12 downto 12));
    hc_29 <= hc_sl(not hc_uns(hc_28));
    hc_26 <= hc_sl(hc_5(13 downto 13));
    hc_27 <= hc_sl(not hc_uns(hc_26));
    hc_24 <= hc_sl(hc_5(14 downto 14));
    hc_25 <= hc_sl(not hc_uns(hc_24));
    hc_22 <= hc_sl(hc_5(15 downto 15));
    hc_23 <= hc_sl(not hc_uns(hc_22));
    hc_20 <= hc_sl(hc_5(16 downto 16));
    hc_21 <= hc_sl(not hc_uns(hc_20));
    hc_18 <= hc_sl(hc_5(17 downto 17));
    hc_19 <= hc_sl(not hc_uns(hc_18));
    hc_16 <= hc_sl(hc_5(18 downto 18));
    hc_17 <= hc_sl(not hc_uns(hc_16));
    hc_14 <= hc_sl(hc_5(19 downto 19));
    hc_15 <= hc_sl(not hc_uns(hc_14));
    hc_12 <= hc_sl(hc_5(20 downto 20));
    hc_13 <= hc_sl(not hc_uns(hc_12));
    hc_10 <= hc_sl(hc_5(21 downto 21));
    hc_11 <= hc_sl(not hc_uns(hc_10));
    hc_8 <= hc_sl(hc_5(22 downto 22));
    hc_9 <= hc_sl(not hc_uns(hc_8));
    hc_5 <= hc_slv(hc_uns(a) - hc_uns(hc_4));
    hc_6 <= hc_sl(hc_5(23 downto 23));
    hc_7 <= hc_sl(not hc_uns(hc_6));
    hc_54 <= hc_7 & hc_9 & hc_11 & hc_13 & hc_15 & hc_17 & hc_19 & hc_21 & hc_23 & hc_25 & hc_27 & hc_29 & hc_31 & hc_33 & hc_35 & hc_37 & hc_39 & hc_41 & hc_43 & hc_45 & hc_47 & hc_49 & hc_51 & hc_53;
    hc_3 <= hc_sl(a(23 downto 23));
    with to_integer(hc_uns(hc_3)) select hc_55 <= 
        a when 0,
        hc_54 when others;
    hc_56 <= hc_sl(hc_55(0 downto 0));
    hc_80 <= hc_56 & hc_57 & hc_58 & hc_59 & hc_60 & hc_61 & hc_62 & hc_63 & hc_64 & hc_65 & hc_66 & hc_67 & hc_68 & hc_69 & hc_70 & hc_71 & hc_72 & hc_73 & hc_74 & hc_75 & hc_76 & hc_77 & hc_78 & hc_79;
    hc_81 <= hc_sl(hc_80(0 downto 0));
    hc_83 <= hc_sl(hc_uns(hc_81) or hc_uns(hc_82));
    hc_87 <= hc_sl(hc_uns(hc_83) or hc_uns(hc_86));
    hc_95 <= hc_sl(hc_uns(hc_87) or hc_uns(hc_94));
    hc_111 <= hc_sl(hc_uns(hc_95) or hc_uns(hc_110));
    hc_127 <= hc_sl(hc_uns(hc_111) or hc_uns(hc_126));
    with to_integer(hc_uns(hc_127)) select hc_176 <= 
        hc_128 when 0,
        hc_175 when others;
    hc_178 <= hc_sl(hc_uns(hc_176) = hc_uns(hc_177));
    with to_integer(hc_uns(hc_178)) select hc_936 <= 
        hc_934 when 0,
        hc_935 when others;

    -- aliases

    -- output assignments
    b <= hc_936;

end architecture;
