library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity int_to_float is
    port (
        a : in std_logic_vector (23 downto 0);
        b : out std_logic_vector (32 downto 0)
    );
end entity;

architecture rtl of int_to_float is

    -- conversion functions
    function hc_uns(a : std_logic)        return unsigned         is variable b : unsigned(0 downto 0); begin b(0) := a; return b; end;
    function hc_uns(a : std_logic_vector) return unsigned         is begin return unsigned(a); end;
    function hc_sgn(a : std_logic)        return signed           is variable b : signed(0 downto 0); begin b(0) := a; return b; end;
    function hc_sgn(a : std_logic_vector) return signed           is begin return signed(a); end;
    function hc_sl (a : std_logic_vector) return std_logic        is begin return a(a'right); end;
    function hc_sl (a : unsigned)         return std_logic        is begin return a(a'right); end;
    function hc_sl (a : signed)           return std_logic        is begin return a(a'right); end;
    function hc_sl (a : boolean)          return std_logic        is begin if a then return '1'; else return '0'; end if; end;
    function hc_slv(a : std_logic_vector) return std_logic_vector is begin return a; end;
    function hc_slv(a : unsigned)         return std_logic_vector is begin return std_logic_vector(a); end;
    function hc_slv(a : signed)           return std_logic_vector is begin return std_logic_vector(a); end;

    -- signal declarations
    signal hc_161 : std_logic;
    constant hc_159 : std_logic_vector (7 downto 0) := "00010111";
    signal hc_160 : std_logic;
    signal hc_162 : std_logic;
    signal hc_157 : std_logic;
    constant hc_155 : std_logic_vector (7 downto 0) := "00010110";
    signal hc_156 : std_logic;
    signal hc_158 : std_logic;
    signal hc_153 : std_logic;
    constant hc_151 : std_logic_vector (7 downto 0) := "00010101";
    signal hc_152 : std_logic;
    signal hc_154 : std_logic;
    signal hc_149 : std_logic;
    constant hc_147 : std_logic_vector (7 downto 0) := "00010100";
    signal hc_148 : std_logic;
    signal hc_150 : std_logic;
    signal hc_145 : std_logic;
    constant hc_143 : std_logic_vector (7 downto 0) := "00010011";
    signal hc_144 : std_logic;
    signal hc_146 : std_logic;
    signal hc_141 : std_logic;
    constant hc_139 : std_logic_vector (7 downto 0) := "00010010";
    signal hc_140 : std_logic;
    signal hc_142 : std_logic;
    signal hc_137 : std_logic;
    constant hc_135 : std_logic_vector (7 downto 0) := "00010001";
    signal hc_136 : std_logic;
    signal hc_138 : std_logic;
    signal hc_133 : std_logic;
    constant hc_131 : std_logic_vector (7 downto 0) := "00010000";
    signal hc_132 : std_logic;
    signal hc_134 : std_logic;
    signal hc_129 : std_logic;
    constant hc_127 : std_logic_vector (7 downto 0) := "00001111";
    signal hc_128 : std_logic;
    signal hc_130 : std_logic;
    signal hc_125 : std_logic;
    constant hc_123 : std_logic_vector (7 downto 0) := "00001110";
    signal hc_124 : std_logic;
    signal hc_126 : std_logic;
    signal hc_121 : std_logic;
    constant hc_119 : std_logic_vector (7 downto 0) := "00001101";
    signal hc_120 : std_logic;
    signal hc_122 : std_logic;
    signal hc_117 : std_logic;
    constant hc_115 : std_logic_vector (7 downto 0) := "00001100";
    signal hc_116 : std_logic;
    signal hc_118 : std_logic;
    signal hc_113 : std_logic;
    constant hc_111 : std_logic_vector (7 downto 0) := "00001011";
    signal hc_112 : std_logic;
    signal hc_114 : std_logic;
    signal hc_109 : std_logic;
    constant hc_107 : std_logic_vector (7 downto 0) := "00001010";
    signal hc_108 : std_logic;
    signal hc_110 : std_logic;
    signal hc_105 : std_logic;
    constant hc_103 : std_logic_vector (7 downto 0) := "00001001";
    signal hc_104 : std_logic;
    signal hc_106 : std_logic;
    signal hc_101 : std_logic;
    constant hc_99 : std_logic_vector (7 downto 0) := "00001000";
    signal hc_100 : std_logic;
    signal hc_102 : std_logic;
    signal hc_97 : std_logic;
    constant hc_95 : std_logic_vector (7 downto 0) := "00000111";
    signal hc_96 : std_logic;
    signal hc_98 : std_logic;
    signal hc_93 : std_logic;
    constant hc_91 : std_logic_vector (7 downto 0) := "00000110";
    signal hc_92 : std_logic;
    signal hc_94 : std_logic;
    signal hc_89 : std_logic;
    constant hc_87 : std_logic_vector (7 downto 0) := "00000101";
    signal hc_88 : std_logic;
    signal hc_90 : std_logic;
    signal hc_85 : std_logic;
    constant hc_83 : std_logic_vector (7 downto 0) := "00000100";
    signal hc_84 : std_logic;
    signal hc_86 : std_logic;
    signal hc_81 : std_logic;
    constant hc_79 : std_logic_vector (7 downto 0) := "00000011";
    signal hc_80 : std_logic;
    signal hc_82 : std_logic;
    signal hc_77 : std_logic;
    constant hc_75 : std_logic_vector (7 downto 0) := "00000010";
    signal hc_76 : std_logic;
    signal hc_78 : std_logic;
    signal hc_73 : std_logic;
    constant hc_71 : std_logic_vector (7 downto 0) := "00000001";
    signal hc_72 : std_logic;
    signal hc_74 : std_logic;
    signal hc_69 : std_logic;
    constant hc_67 : std_logic_vector (7 downto 0) := "00000000";
    signal hc_68 : std_logic;
    signal hc_70 : std_logic;
    signal hc_66 : std_logic;
    signal hc_65 : std_logic;
    signal hc_64 : std_logic;
    signal hc_63 : std_logic;
    signal hc_62 : std_logic;
    signal hc_61 : std_logic;
    signal hc_60 : std_logic;
    constant hc_54 : std_logic_vector (23 downto 0) := "000000000000000000000001";
    signal hc_51 : std_logic;
    signal hc_52 : std_logic;
    signal hc_49 : std_logic;
    signal hc_50 : std_logic;
    signal hc_47 : std_logic;
    signal hc_48 : std_logic;
    signal hc_45 : std_logic;
    signal hc_46 : std_logic;
    signal hc_43 : std_logic;
    signal hc_44 : std_logic;
    signal hc_41 : std_logic;
    signal hc_42 : std_logic;
    signal hc_39 : std_logic;
    signal hc_40 : std_logic;
    signal hc_37 : std_logic;
    signal hc_38 : std_logic;
    signal hc_35 : std_logic;
    signal hc_36 : std_logic;
    signal hc_33 : std_logic;
    signal hc_34 : std_logic;
    signal hc_31 : std_logic;
    signal hc_32 : std_logic;
    signal hc_29 : std_logic;
    signal hc_30 : std_logic;
    signal hc_27 : std_logic;
    signal hc_28 : std_logic;
    signal hc_25 : std_logic;
    signal hc_26 : std_logic;
    signal hc_23 : std_logic;
    signal hc_24 : std_logic;
    signal hc_21 : std_logic;
    signal hc_22 : std_logic;
    signal hc_19 : std_logic;
    signal hc_20 : std_logic;
    signal hc_17 : std_logic;
    signal hc_18 : std_logic;
    signal hc_15 : std_logic;
    signal hc_16 : std_logic;
    signal hc_13 : std_logic;
    signal hc_14 : std_logic;
    signal hc_11 : std_logic;
    signal hc_12 : std_logic;
    signal hc_9 : std_logic;
    signal hc_10 : std_logic;
    signal hc_7 : std_logic;
    signal hc_8 : std_logic;
    signal hc_5 : std_logic;
    signal hc_6 : std_logic;
    signal hc_53 : std_logic_vector (23 downto 0);
    signal hc_55 : std_logic_vector (23 downto 0);
    signal hc_56 : std_logic_vector (23 downto 0);
    signal hc_58 : std_logic_vector (7 downto 0);
    signal hc_1 : std_logic_vector (7 downto 0);
    signal hc_59 : std_logic;
    signal hc_4 : std_logic;
    signal hc_163 : std_logic_vector (32 downto 0);

begin

    -- logic
    hc_161 <= hc_sl(hc_56(0 downto 0));
    hc_160 <= hc_sl(hc_uns(hc_159) < hc_uns(hc_1));
    hc_162 <= hc_sl(hc_uns(hc_160) and hc_uns(hc_161));
    hc_157 <= hc_sl(hc_56(1 downto 1));
    hc_156 <= hc_sl(hc_uns(hc_155) < hc_uns(hc_1));
    hc_158 <= hc_sl(hc_uns(hc_156) and hc_uns(hc_157));
    hc_153 <= hc_sl(hc_56(2 downto 2));
    hc_152 <= hc_sl(hc_uns(hc_151) < hc_uns(hc_1));
    hc_154 <= hc_sl(hc_uns(hc_152) and hc_uns(hc_153));
    hc_149 <= hc_sl(hc_56(3 downto 3));
    hc_148 <= hc_sl(hc_uns(hc_147) < hc_uns(hc_1));
    hc_150 <= hc_sl(hc_uns(hc_148) and hc_uns(hc_149));
    hc_145 <= hc_sl(hc_56(4 downto 4));
    hc_144 <= hc_sl(hc_uns(hc_143) < hc_uns(hc_1));
    hc_146 <= hc_sl(hc_uns(hc_144) and hc_uns(hc_145));
    hc_141 <= hc_sl(hc_56(5 downto 5));
    hc_140 <= hc_sl(hc_uns(hc_139) < hc_uns(hc_1));
    hc_142 <= hc_sl(hc_uns(hc_140) and hc_uns(hc_141));
    hc_137 <= hc_sl(hc_56(6 downto 6));
    hc_136 <= hc_sl(hc_uns(hc_135) < hc_uns(hc_1));
    hc_138 <= hc_sl(hc_uns(hc_136) and hc_uns(hc_137));
    hc_133 <= hc_sl(hc_56(7 downto 7));
    hc_132 <= hc_sl(hc_uns(hc_131) < hc_uns(hc_1));
    hc_134 <= hc_sl(hc_uns(hc_132) and hc_uns(hc_133));
    hc_129 <= hc_sl(hc_56(8 downto 8));
    hc_128 <= hc_sl(hc_uns(hc_127) < hc_uns(hc_1));
    hc_130 <= hc_sl(hc_uns(hc_128) and hc_uns(hc_129));
    hc_125 <= hc_sl(hc_56(9 downto 9));
    hc_124 <= hc_sl(hc_uns(hc_123) < hc_uns(hc_1));
    hc_126 <= hc_sl(hc_uns(hc_124) and hc_uns(hc_125));
    hc_121 <= hc_sl(hc_56(10 downto 10));
    hc_120 <= hc_sl(hc_uns(hc_119) < hc_uns(hc_1));
    hc_122 <= hc_sl(hc_uns(hc_120) and hc_uns(hc_121));
    hc_117 <= hc_sl(hc_56(11 downto 11));
    hc_116 <= hc_sl(hc_uns(hc_115) < hc_uns(hc_1));
    hc_118 <= hc_sl(hc_uns(hc_116) and hc_uns(hc_117));
    hc_113 <= hc_sl(hc_56(12 downto 12));
    hc_112 <= hc_sl(hc_uns(hc_111) < hc_uns(hc_1));
    hc_114 <= hc_sl(hc_uns(hc_112) and hc_uns(hc_113));
    hc_109 <= hc_sl(hc_56(13 downto 13));
    hc_108 <= hc_sl(hc_uns(hc_107) < hc_uns(hc_1));
    hc_110 <= hc_sl(hc_uns(hc_108) and hc_uns(hc_109));
    hc_105 <= hc_sl(hc_56(14 downto 14));
    hc_104 <= hc_sl(hc_uns(hc_103) < hc_uns(hc_1));
    hc_106 <= hc_sl(hc_uns(hc_104) and hc_uns(hc_105));
    hc_101 <= hc_sl(hc_56(15 downto 15));
    hc_100 <= hc_sl(hc_uns(hc_99) < hc_uns(hc_1));
    hc_102 <= hc_sl(hc_uns(hc_100) and hc_uns(hc_101));
    hc_97 <= hc_sl(hc_56(16 downto 16));
    hc_96 <= hc_sl(hc_uns(hc_95) < hc_uns(hc_1));
    hc_98 <= hc_sl(hc_uns(hc_96) and hc_uns(hc_97));
    hc_93 <= hc_sl(hc_56(17 downto 17));
    hc_92 <= hc_sl(hc_uns(hc_91) < hc_uns(hc_1));
    hc_94 <= hc_sl(hc_uns(hc_92) and hc_uns(hc_93));
    hc_89 <= hc_sl(hc_56(18 downto 18));
    hc_88 <= hc_sl(hc_uns(hc_87) < hc_uns(hc_1));
    hc_90 <= hc_sl(hc_uns(hc_88) and hc_uns(hc_89));
    hc_85 <= hc_sl(hc_56(19 downto 19));
    hc_84 <= hc_sl(hc_uns(hc_83) < hc_uns(hc_1));
    hc_86 <= hc_sl(hc_uns(hc_84) and hc_uns(hc_85));
    hc_81 <= hc_sl(hc_56(20 downto 20));
    hc_80 <= hc_sl(hc_uns(hc_79) < hc_uns(hc_1));
    hc_82 <= hc_sl(hc_uns(hc_80) and hc_uns(hc_81));
    hc_77 <= hc_sl(hc_56(21 downto 21));
    hc_76 <= hc_sl(hc_uns(hc_75) < hc_uns(hc_1));
    hc_78 <= hc_sl(hc_uns(hc_76) and hc_uns(hc_77));
    hc_73 <= hc_sl(hc_56(22 downto 22));
    hc_72 <= hc_sl(hc_uns(hc_71) < hc_uns(hc_1));
    hc_74 <= hc_sl(hc_uns(hc_72) and hc_uns(hc_73));
    hc_69 <= hc_sl(hc_56(23 downto 23));
    hc_68 <= hc_sl(hc_uns(hc_67) < hc_uns(hc_1));
    hc_70 <= hc_sl(hc_uns(hc_68) and hc_uns(hc_69));
    hc_66 <= hc_sl(hc_1(0 downto 0));
    hc_65 <= hc_sl(hc_1(1 downto 1));
    hc_64 <= hc_sl(hc_1(2 downto 2));
    hc_63 <= hc_sl(hc_1(3 downto 3));
    hc_62 <= hc_sl(hc_1(4 downto 4));
    hc_61 <= hc_sl(hc_1(5 downto 5));
    hc_60 <= hc_sl(hc_1(6 downto 6));
    hc_51 <= hc_sl(a(0 downto 0));
    hc_52 <= hc_sl(not hc_uns(hc_51));
    hc_49 <= hc_sl(a(1 downto 1));
    hc_50 <= hc_sl(not hc_uns(hc_49));
    hc_47 <= hc_sl(a(2 downto 2));
    hc_48 <= hc_sl(not hc_uns(hc_47));
    hc_45 <= hc_sl(a(3 downto 3));
    hc_46 <= hc_sl(not hc_uns(hc_45));
    hc_43 <= hc_sl(a(4 downto 4));
    hc_44 <= hc_sl(not hc_uns(hc_43));
    hc_41 <= hc_sl(a(5 downto 5));
    hc_42 <= hc_sl(not hc_uns(hc_41));
    hc_39 <= hc_sl(a(6 downto 6));
    hc_40 <= hc_sl(not hc_uns(hc_39));
    hc_37 <= hc_sl(a(7 downto 7));
    hc_38 <= hc_sl(not hc_uns(hc_37));
    hc_35 <= hc_sl(a(8 downto 8));
    hc_36 <= hc_sl(not hc_uns(hc_35));
    hc_33 <= hc_sl(a(9 downto 9));
    hc_34 <= hc_sl(not hc_uns(hc_33));
    hc_31 <= hc_sl(a(10 downto 10));
    hc_32 <= hc_sl(not hc_uns(hc_31));
    hc_29 <= hc_sl(a(11 downto 11));
    hc_30 <= hc_sl(not hc_uns(hc_29));
    hc_27 <= hc_sl(a(12 downto 12));
    hc_28 <= hc_sl(not hc_uns(hc_27));
    hc_25 <= hc_sl(a(13 downto 13));
    hc_26 <= hc_sl(not hc_uns(hc_25));
    hc_23 <= hc_sl(a(14 downto 14));
    hc_24 <= hc_sl(not hc_uns(hc_23));
    hc_21 <= hc_sl(a(15 downto 15));
    hc_22 <= hc_sl(not hc_uns(hc_21));
    hc_19 <= hc_sl(a(16 downto 16));
    hc_20 <= hc_sl(not hc_uns(hc_19));
    hc_17 <= hc_sl(a(17 downto 17));
    hc_18 <= hc_sl(not hc_uns(hc_17));
    hc_15 <= hc_sl(a(18 downto 18));
    hc_16 <= hc_sl(not hc_uns(hc_15));
    hc_13 <= hc_sl(a(19 downto 19));
    hc_14 <= hc_sl(not hc_uns(hc_13));
    hc_11 <= hc_sl(a(20 downto 20));
    hc_12 <= hc_sl(not hc_uns(hc_11));
    hc_9 <= hc_sl(a(21 downto 21));
    hc_10 <= hc_sl(not hc_uns(hc_9));
    hc_7 <= hc_sl(a(22 downto 22));
    hc_8 <= hc_sl(not hc_uns(hc_7));
    hc_5 <= hc_sl(a(23 downto 23));
    hc_6 <= hc_sl(not hc_uns(hc_5));
    hc_53 <= hc_6 & hc_8 & hc_10 & hc_12 & hc_14 & hc_16 & hc_18 & hc_20 & hc_22 & hc_24 & hc_26 & hc_28 & hc_30 & hc_32 & hc_34 & hc_36 & hc_38 & hc_40 & hc_42 & hc_44 & hc_46 & hc_48 & hc_50 & hc_52;
    hc_55 <= hc_slv(hc_uns(hc_53) + hc_uns(hc_54));
    with to_integer(hc_uns(hc_4)) select hc_56 <= 
        a when 0,
        hc_55 when others;
    the_priorityEncoder: entity work.priorityEncoder (rtl)
        port map ( a => hc_56, priority => hc_58(7 downto 0) );
    hc_1 <= hc_58;
    hc_59 <= hc_sl(hc_1(7 downto 7));
    hc_4 <= hc_sl(a(23 downto 23));
    hc_163 <= hc_4 & hc_59 & hc_60 & hc_61 & hc_62 & hc_63 & hc_64 & hc_65 & hc_66 & hc_70 & hc_74 & hc_78 & hc_82 & hc_86 & hc_90 & hc_94 & hc_98 & hc_102 & hc_106 & hc_110 & hc_114 & hc_118 & hc_122 & hc_126 & hc_130 & hc_134 & hc_138 & hc_142 & hc_146 & hc_150 & hc_154 & hc_158 & hc_162;

    -- aliases

    -- output assignments
    b <= hc_163;

end architecture;
